PK   �[^Wu����  ��     cirkitFile.json�[��6��J�}��.�۶���&�,���![TG�c�j�m����|["�c�3N��C�1υ"?���˨)>��t�j���m���rt��x�X4�����t<z����j�kS<=������O6��>>��v��jc�a�"�x�9Ku���y2��r>���l���><��VgN=�<cE%
���,��$�R$����\�\�S�F��:Ÿ�F�8u�S�8u�S�p�y��M�jY�XaL"��&E>���X�f���8b0���(�CR��G�ΐ�3$�Lc�N���`\��C5���9rj�H�9�z���#��
3��5�"'	��%x���QC���X�g��v�5ױL:9"\�29`F��,P�#�A�ģ#H=a�F<��m�%l�����,��ZM�V�Y&���d681�c��<��1H=������� �x. R��0X��#i?� ��� L�ޙ����!�;�������IEa��h�<�U��t��D��$��t��j&+��Y�F��0ױxr���m|�kT����~���\'��"q*�ʹJ
k�TΤ(�D6xl�	r�k��b��ౄ�rc|�v�2�͠2vh���\#�S�ʻ�K,�o�\,�s�@��9�\,�s�D��9K$��J$ɟD�'��I$ɟB��)$
ɟ�.���)$
ɟB��i$ɟF����p0;����m��׍x��ϱm]���:��	\Fa\��r���Zb\�<8p� �����^�|�X5��JFK�?#��%ފ�L �po��l��� y"IbE�X�$V����J�Z�r^0u-�nNI3�1�h� �1C�/����hff!�fh f9�N�9Ŝ�bNC1����-7�ř����DbNC1χ��+l(�C�S8?�@�98߼����m�����b A]6�����ఆ��X��� (�#������
�� ����+��fhί�oPD=���+�+>Wg���R���P�ϯ��I&���
|TNQ�|(�`��F�ߩ,4���ł�bA�M,4�X,hb���Œ&K�%QFLC���X�P,i(�4K�Ŋ�bEC���X-�h(V4+�Ŋ�bMC���X�P�)�~XaC	$�P�|]���u\�@O}�?� ��
z{x��c��u���cեݬ�b�<V�[�$V�IbE�X�$V����JNC�4�2|��`FC0�A��0�h f4s�9Q����P�i(�4s�9Ŝ�b>H1�Xoe�a�*�� ��cU���v��д�����k�*����PG/����X������X������X� ��P<�_��U	��P<�_��U	��P<�_��U	��P,h(4�T��bAC���X�P,h(4�%Œ�bIC�$ʈi(�4K�%Œ�bIC���X�P�h(V4+��Ŋ�bEC���X�P�i(�4k�� ��cU��������e���Ǫx+�O>V�[�:v��}���:���Gw\�G���>O��ܖ�z9]5�mFw0_Ë:yc�7uކq�Q�Ϙ���r���
�����&����]��������a�[��HP���V�z�H8���`�:N�g8���s����Pۣר��^�L�������#��i�kt60O��.4^��_tEC��.\LA^�{xدM�q��-N�eZ�|p�t�'�~����5�ȥ�����fas�
���_�
�t��·ZnxB�;�/�
�_�q��'�#�A����`�*`����*�7vq�o�����-���
 ��g+p��;��5�إ�H�.�cQb��\�p�N@� "���8o������F��l�|�<45�d����6(>�GESn���.���UUm�����^�b��~z�'�T��/�+Ø��H}���H}��ϐ�y�;1;l��=Ԟ!��ϱ��2,��h{E��)�]Lӷ���e��Hd9�S��c9�XN۫(*4�6�rlpm�t�(����۱Y�o���!�
0,v��æ�`X�������j�g�a�z�tg�,�`�������?3!����`�<�8�o��`!<�8����`9<��o����s���n'����uf$��"y�Jo�rתg��O�Q_ʲP�Ȳ0�!ifK]�wd�7�1LR+̀��-��[`��n���%6pKl��X0%6��X%�D�%QbI�X%�D�%QaITX�D�^QaITX�D�%QaI�X5�D�%Q�!|����a����;D�1�Wna�%��-,�_�혋d��۸s�D|-�c.�Ɓ��v�IQ��L]��Mg��pB�@�o����V����������}^�sa�P�e۾m������ږb^�y�5���m���F��I�N ���0��ͷd�_i����u��������^Cx�5��^�}�Xz�5�א�x�5�א^Cz�5��P^Cy�5T��^Cy�5��P^C{�5���m�Bb�K�:es����Ga��e�%���IYZ��Ҧ6���z�H?��~�#����f;B�v��t��'�os���Ꮸ��{�� Q���i�2�{��z�67�*�߰�T}{��߃��Bu�����w���M��A_��g�����>t?FT{E��Z�+s�����Q����� Q�u�~^��mn���~DmЗr�+Dm�oi��`k��B�bf>�� ��ٮ�xw��+b�"�+��"�+�"�+R�"�+��"�+��"�+2��lW����]Q�+b��`��`���۷�7�7��?6�?7۷�7۷�����b���[��U��[��j����?m�P�ɓ��U"�2�,Y��E)SY��;+S>�w�q��$?�c�����V�v���p�0~�G�.�g_ڏ�5�'۬k�W������u�Z:������Z��5��L�Ts�,z�t��Q��|n*Ѥ�餓,˙�p�T�Ȅ�m�n%�.��h=>���U���h�yr��f�����ࢨ��X�0�����`�K�q�<.��%쨄�f"��ZJ2+�Q�Q�Ic:,��l�J��KS�0�%�D���vTh�}I���%��ڗ��j_�o�}I���%��ڕ�ʗ<���V�߯7e���6�[�؄M�΁�3������A�$��M���Ѻ,>��}�x��Xl�O����}x�,k7BG�Ϗ��o��;ˣ��X<[W�l�_��z������M�X7��.�!��Xn�b��4�k�U8;��S����͒�*�𡅜��Fi���L�L����
Q��d��]�+��$��yɜ�����hO�8���J{��lY������ZF�8�.���I��nb�!�"��Jնp,ro�u�R��S�N@ߚ���E�l����������iՙ�Z��	VZ��2f�dy1K�,7��r�dL�J�Y%̼�h�0i�� 1����?w�L��U梴�5�gFOR��L��P�\uR���� �,`�g�Z��BNb!�L���BNb�9�AR���G��
xH<*P��R����ǀT�#=c@*�1 ��S)�]��D�gH��HAj�"�h�ӷ�kʓ�T�������Ӱ�me�o뚂�ڗ
ԗ
��ǀT���Tȣ�<c@*�/�A�ؗ
y�K�%�c_*8.A�U�R!�}��ǴS/v���f�,�ikh�ܖ���mI�ګ�<k�w�?��:�%���;�K��N��$[���B�R&v6���ʊ�ԙM29+�L+f�m��lt �VY��<m3Q����)��;_p��>:�g�f/��+�7��ͣm��r�Z��To~x��gz <�ES��8�t����蓝3�!v��O�Gբ~�~�������^?�;�n�\mf���_��fY~�*��R/��ʼ4��-�U{7�����}*�Or��:�ag����x�_J�j���|���r�����
Fy:h-j�j߯6n 4o~���U�;p�	g*�8�\I#��5f��LK����t�S��k9�I!�<)�L&�f"Ѭ*
��;O����2<|_=^���w	c��+�.��>Un&Lfi��$��v��1�us�y!�MĬ�I��2>�r�S��EV��$N��.d��u68�����\�J��m�0����ᆄ�K\ Z�{P&�2(1i��s�O��,�R�^=��p+9�I���ۮw��011���#������[H�Kp���G[���E�Fj���%�߻����/{�G[~w8�z�����_j��?�����ڗ�Q�k[�Gw�~���v?�;������˶����ZkvY��{_�5��ߓ�����zO��e@��������~��V�|��v`>�O�>���GK��ʼ�8(&UPL	s���a��m�3b_�G_y���;�,)E)E�����"vE\��!D�߻b)���l�/��+Ō�g�쉅�L����ɜIN�dNJ$����~�y*��H$��
��adW�$,^,�BD�ǟa��[o�QR�!)���&eR\7�f4�v�D�����w@����.k��L��b�b�g &��C�� �K�wq�LATv�b��R"���u��1A)}�'�~=�a�6��5������]ʣ��cW,��RRE��ҠR|�ǾP����y̩yT�<�k�h|�鰘�B*�>�������hb	�k��NJ� ٯ��k:b܄��R�t�3�$:��b٣�L��hi$�����}��R%J�E=�Tl���&�BbcO� w��W$���0^P5���Oߏ�
���y��ڷ|��|WN��}g�'�r������;{|��<��}��˫�2�.�ݽ%�
��ԍl���և'�_�wN^�	�a�r�g�.��]N�5E���&;]�6���	��0�sC�崑}W=\��p�vڛ !�AG��vU���/��.�Y�_wdw���Ԅ��N.�����]]0�a_�@��$pԍ�ϯ;|���	�N�C�^%�þv���%q��vI��d�C�b�ݿW/o����m�b�<��<�?���b�)߭>����}M����PK   �[^W���[�� f� /   images/8959c7fa-44e8-4699-8891-15a891fa383e.png�eT\]�.
4���i��-�4�n���%x������	���������q�;���W��Y���̪U�V��p��RH�x�```H2���``��``B��q�g���SUMge��������	��7{wS00��/:�}$�������E2��D]~�
�����p/7A��;x�Z͍�2Mkʩ~K��ʜv�Kzϝ[�0��	�q���в;z��%J�bɉ�]�*���a�����/���hu�jY`oJ��̩��x]�VW�������|I�0q��G�;;�I���V��0�3��rM�}��_Al�5�F�56^1���e��X���제c�W��D�%��S��_vX��;^@�O�`@_�P��md�wYB���S��|o��3�^&�TO��֐�|π����+�����s<��"�v���Z����X�P�<�y�MQ"K��'@�!�0r:������C�^^�WN�1�v,��蓬}��\af�6�7�i��ɏ��{ �9~ux�v���D�L��wH�dp��(7���GS���n-w��)W�,�V|�U���:���BQF)����JW�V�F= �q�A���O�*ZɊÃ�ݲ����\"�E��OpH��o���KX��1ǟ�c������]t��IL�)x*_�e"i����,&<�֟�NZ�u����{���~�.ɭ����Wd&U��mUmM���//�o��q�!��a���
�Fv6L c;C&w{�����=���ę�����V�좭����X�L�C�`/fbn!��h���Y���ʈǘLH�ߝ����D�ncm���.@�.���bf2�T���4�H��MHؙؙ�����d��$��Ʀ�����1 3wv��efvsscrcc�s4cf���a�2��2~h0:}�u�3�:���������������-��1����Y���c�����^A�?�m����`v�3�0�ml���'g	W���3�T?�3�������������3��CH�((�7��,l��1�c9�����?��]���16b6�6�� u�`c�o���������gq����ϖ�����x��\��ʈ��]/�����1�??���\��윌 N�	#�	;#���1#�1��	Д��ߠdl��A�F&�>$L8܆<� 6N.F�����ѐ���d���2arp������GT���}U��?����L�8@l�\,&��\܌��� FSSvvSc.n���^^%2V&�I��AΦv�6d
 #E���Q��1Qq��'7'7������_J�&�N�����/*c#^�H�G�X؀�L��m����{]�Z�a����X����b�& g;GU;;k���$!�sZ�c?��A� g�6 +/������������M�����������C��//K[8}��G��-�b��ѿ������+xAF�2�	�jbL�ߦ��A�f&����-�������cld�h�j�������N#FnnC �Ј��Cw�3uv9���}���WA���Hh�u	i�������|�n�������?,f�w����oN��¿���ً�?��G6d��t�N������!���!���!���_���WCeb�Q�}�K�&��������78X�w�!�����!</�������PNJ���+��81c_F\D�}��"�xQ�	�� ,j�ۯ�<�:�y�R�R��c�F���j�eh#���]�-�I���oW�~�ey��"u�!��D�&Z)�r�)���u��l���n$N�]��J����SU��ݸ�xy�ǜ�v���_�y���ťM�}~�#_l��8�R�jj�_��m�v�~�-�9�C(����z��|uN�6k�m#���d,�s���j����*���Ѩ�9B���mkѰ&�BG�W���Z�
,'ktz�����J�0I�dAA����Ư�ʯ�t�N�-�t��T�0�"$�CW7����xݔ�0��8(�{Yg����=i�Ծ��b�%����'��^�`1/��z�>�K\�K���?o�O��iW�OZsr����C0�����i{m&^x�f�'Ӈt�C��F���x��ਃ�@oN�1��F�܎_����/5���*���=��m�|L���q�J��Q�H,���:�������ܛ���acXw�u�I�+Y�j�H���쥏�	�k��I�A�u
`7�['�_�lio;�
�&��v�Z1�{zz��COs\k
�p���i����'=�L��G�v��1�e�R�}��J��e������>��Z���� <Ld�՚S_E%p��~,����}�G	��bnd���~�A�+OL\�p�ٙ�B��5ذ�GUy]��R��@�8
�����t5���ϛ�|��n���m`� �.@������rѝ�3(zv��6�<�>�N��%Ҡ�"%�~8�+^��e�4$�^���5,m2����`%9���.9�w)'�4wJ�n�(�FJ�`O�%ϗ��f�Ρt�B��p��:�n���ZY��O9&����#Ƶ���Ĺ�X��VVVW�z��a��±J��R]V�DAcj���d�x^��W�pcl,�܉�*�[���4����m�U���{Т'(��Y�i����敒/'K7�%3�U~�:}m��O��!n��=?��$g�
3�6 3��[�]r/�F%a������)v��h�XC�Z˞
�`�rĚz��OY���f�_��[r^�\{�Z�bts�i���<��J��U�ܪ�Hɤ��A�2��l�
�g�5��X�;C,��C+��؋�-�:Q�u�AN�Iμ�|����R��v
���i饿��rqq�0�Gܶ ����|4��%Uě`a���s�� ��D|kf;��F����L��~�ǻ�،Ք��#�C�O�aE��	_�M�H%bKk3���ĂҬ�v�e����{юt�yްځ1ީN���HOj3�*��j1�l��S�,z8��>O���wvp2b�k��W�2	�t�p2X�h���qJ@tĐ��=�q�������#�bZ8��/�#�Â.-A��^�*[%Lj���Y%§�����L��͹�02d�E����������Z�md��ߠ�:kE�"<b>��xe�	�URw�ʅ��Mʇ�E��]���N_�a�@��G��s8�{�jr7A~�@���.��m�4���-zü�(���f�4^�p퐺�8D�d��x2�R�d9�]��Ŕh��D�r������{�|����t��?�)���5f�����p�����i�
l���?��I��w�Kk-�~)ko�o�S�����f�O�G�8%�MQ%,~LI5���r���W(e�<��0#K�+��A	���ot��+f�b�''v>Mؽ�����H�ytm��3��=~�%~��q���XC�q|�y�f|©m�kе�����W����Z􎴋Ji�k~q8>p/R�(f��'������p������I� ��\�`�}�����u�/�Eש�*xM[{�/	�	�h{���-/�e$~���<���6%��L�wi�C!N�uv3Qp/+��Z-�z�Eu(T���~t) Q�1(�9,?h�ޮ������R��F:u�Le��z5�Rs�ȣ`L���ծ��"�m�v�hJ:2��Q��Ո=XO��u���tt�
vք[��T�q\�6�`I%��IB��j�<�k��̵�v<7�;���F�l?捲����o4)�t�ɿ�<6�jUsKD�Ӑ�G~Mm;r�pnĜ���!PF摱�r�~dxLlj@S�`.C��L�����,���`�������I ������_w�Zg�
_�,��S@�k�*�so�ɑ_h�w�[T5 ����l��bch����c���4r̈���Iq��'�:~�>���&�2�5Q�?��"��l��"��~��� �m��U�/��7�r���U6ʌ<�~(ڂpKD��ᓈ5\D��=bW��d �����[���v���F�;�=�.��
�k�G�{Q�nTz �!�yE��2}��.i���x�����}�1��I��Z
�1=�]l\~o��������4sl �٘�<�]��i�V~M�-��q��,���nk�N�����v�r�h�q>J�s���*��G��:នS�fS�p���^�pg��D�o}9��48zhe��"���t��=)3��_����8�&�F��ؒL7������d�*��ـ
*�����q��'���_�F��`(a�+5-��p},��sl���\�t��7��N���`�;MƄ��Y�yG"�O����?��**���L�es7{G�1�K$�<�s?O��C&�{��{E�{M}�~�a�60 �[op���݇:me'y��y���:�׆�����2�A<�ﺦ��}�MI)���7�N�Y0�����G�5o�%��vX������P���i{���?�KY���-�'Il�@qU2��-3�J�6.�6栗[���`��
�&<�%���Қ����S:Ծ��&�\��v	QH�%�!��ɉ�G�k�-$�!�)���jqppК���*]ґ���1�M%]���$Q`r.x�:��㠻�,������#�=��A�4 �)C��;����B98��w!@\PS5��4�S�X%���ۢ�v7���vr����I#�5�MЖGؤ���JKxT� ��eJ�_�J%�_��W��[K�^cä�VM5V�A�H	����Q��.������`��V �̱XfTW���Gu�3m@�@P�#��U���%������YB�@BsI����y0&?gh��E��~|���uh�sƽ��3C�>�	2َ�:�F^�>S|�z�2I�b8�5��	`�v�/�)e'�
2�A�u]�>"�M-9����n+�?���ej>{�ఌ���Qžq.�,���],�Js����.����q�3��Շ��0�`�~=�go%��mG�F�YMHO��u��0#��>�&�WͶ � ޮu�~�Pʢ��w2ЩE��J5�ךA1O;��x�=���E�wb�6@:x�V�I��p��qÖ�C������-w�ߘmbm�kx��K�zӌ>����xf�=/�#l��+���:(�"�)n'
�i�&Yg�
t���2[W����c����%��MP+�q���=X"�#g�����=�ֆ�}��1�]��v���v�$U�S	�y��y4] �p�'?�?6k�$V���ܹ���?���͸a��amUoZ�z%,� �X�����x���P�����E�R7�؅���YR��_�vP������ѕ�X1�����3�}�B���T��l]�h��^�V�Z�


Y<N�3���*���ET�������\�<NkSSS\�W�V�LTd����-L����<=ͥ��������tաk�_Tl4w<c�-��M�2"x��Q��.p�P�g����烓���111!!!���[���[/����� ���H�+�9��<��%���܉�{8�mX�N8�g�\kv~~~q��lR/�GM�$� 4 ���c@�ͤ��vNE�[9"�h'&��l��ߜd�W�B!?�����	�G�?��g��xmw�=�A�+[ �*�L�b�]��$�a<�\�X;8(BW6��������\-��k�V�G�&-)%E
o@oh�#D����讴j�1�rmGnpjs3�� }������D۰��T,���;W���?��^��j�
р�����$�xY`�J��zE[L]����-���uaYZ~Ӧ�PP�������7g�F�8���ZD��rr`�G����6ըUx0��P�N��Ƨk�M^Llf�Z�{��.K�i�+�ۣ=�)��x@d*,����c@���Ԧ����9����}RHy��n髕SލY��a	MA���q����k[cqq�.-n�􋼥�5�� ���|߲f�$_���=��T%�%��zĀy�$2nFFƊ��
F��Զ��@"�-D~(��d}� DQ5� �@�26������]�Z����N.v�ҋ3�6��V$�uo�	�i����(��O���,GNi\�(�{��^�'����*z�63�R�R|��`љ�F���I W���d4��Q��ں�d�W���IH�`x{\cބi�!�����sC"�y��c(��(4n�Hy����1w��`\��ID�,x���'��wu����U��M#
�G�Y�AqP��k�m�I������0܎<�rs)���]o5�Di�4�T�9�N�D�0��sk��i�HX}fك<�	,�1�8�y� hFb�r��F�)�� �|��d�s�o�	�{D'�靆4���PyZAג!��f9�*(���.d�f�ӝ��wؒ;ؙQ1]Um$�9XXFH4��V0g�Jz�z<�7�O�/P�M+\������J�����t��u9]t<��HG{>��N�!�"����Opb�:D師��X4d��n�dā2dy���o$�ɮ�̠��H�����f��f�E��(󟧜������=��� ӃT$�s���<E\_9�nb��!���L�D�C��g��8�x��~�9�i���j�7�6.w� ��~��Ov�DV�3�C鈀$L��6��ƉL.�y4��R�@��Xn߫߶����#�]{��n���.���/����Z�ޫ
X�Z����ew~P �"#��M��,�?����(H!���FZ�D�����O��R�i�:�t�6��#�p G��
�."��No>T�-���ӫ)�~����T殛_|i�s|���j3M�OjK+�~�	�0�Hj�$;�}͊2Kals=�5�����H#�l;FA�| ��$����29�S�>��$+��q�g"a榲�g����nZw]����Y�Cd�	�)4A4��!3,(b{|Zб��|��a�I��	@D1qU�Wt��:�ٺ	�z\��?�
L_nu�OAtJfĲ��i�դ;�5ҭS���)�=��<_6�p'aS�2��A�o!A���w�{=�Q��[��(3
n�h��� ���פ5���B!�eW���-���X)�2>�f���7 ��YPGX'CtQ�ǹ�h��Hz_a�#���?]|m�ߞ����){�b�9��1����[Q���CGY�q�,㾙���ՙ׺��~� ")�xyx�m䂢�JTnn|z��zɧ
N(���_��Y���ek5ǐyQqD!�SU�G�ՠ٢h`BL��	-�96�́�X�Aa�ӝسٌ��ƨ���tXn�0% �5��>�lN�=����,A�БӲ�˯h|N1�>N+k��]*�%�1���ݪ�{��C��'�qRM�e]^�)��\Ce�Jl��WQԒ�Eݪ� VOͮ���TH�%2s(�af��Kj�$��ꨆ0�y"[>�������9W�c�F�Y��g.`�J)�E۳�M�� ǚPt~���λۤ�1��4��G�?�bt�,��j�j�:���Ln@��S����Z�����W����x�&���Ͼ6�v�@�ϸ��*�Z{!(�wXsE���聐!����2��f��Aj�?��P�9��3���tD}绽�8�L�#�~1W���R%������k����~�ğ���3�)XT�,`q����۸���5ޕ�9ۛ7�ۄcX�8oq?w��h$jm��C�zg���D6_�9�2zYz��A�:H�{	j�r�k��Vp����������R+�Za��B�"?7OI
����J���އ"�Y!*�����!���g��-G�]k�>Y>؉6����1MtCx��R*���o-��n͉~���F�I>8��j���'�۸Pmn�!���eꇭ��Z��G��~g �/܈��?��x�'�;n�/|����i�e,��9���?D�i9"a#Ke���m�s��p�HBq��N|�{�c�S/��'��&���zY݄&񃝕M3��V�0��\ \̜�#{���w��z���/}I�,�)��o��Nֳ�~ً �����;����5l��#�G=�s/��3-�@*�P:00�u�$�\Nd[�3-6��y7��uWa�����^U���=8�Z�{Q:j���?,�'|�ב3�:iĸ�&��x��9ETY^G�O�IQ��?�A2(Ha ����C(!6V8�?���(��4��m��a�ͨFx��>"f�6��y�<QȟL�N8����9�W:c�r��u�{�&4�ߢy�l� y�%xa���eq]>W�c(EpAC|*M��׬�?����5Sl��>�xDamF��n�<kvȹ�?��R��JM��T,}W�W-��l������_����"��.&;<���}�.�e�ʯ��%����l�	��*+I��Ǆ�L^���D�y���Z1�K����:����t۾���2��i��a�jv�AK���vbCC�OZN_�����2!�������䥰v�(a4p}K�旆T��h;/����	�n
�[nk���i�w�'�mXT���J��O=�0T{��}���6�h�!���j�,|�=���{%M�^we��Ɗs8�P��h�Se�,Cҗ�ܕ���Vk�jf���Z����Sek���"�-^k?}�<���c�R���y�f~�����8 +@�7�z�<����d<�vⅮ j���V��C� I��vpb�(���h�A-ETu<�`22�O� ��sw��60Rs��	�F��i���*937�9?��Bp������)����E�C�է�/�������n&ܨ(�50^*
��x�|��� ��;=B�Pm�H49���5-,�ũU1��ז]�+�mi���T�8nrY�-j��-�ҼHF�NmE�Y�k�T�sArߣ�T25m����H��<�e��|}�x��ň��zb�H���"���u�0�`�ֆ�'��攐4����e��X��aE~p��YsX�U�?���tϾ��`��g������["�"���e�69N4؟ɕ�������� ���X��-�k��ʈ�P�s�uކ�<���zIإ�eV�mp=# l�d�.����a�!ΗJD�eZ�-i^�n�a����XK|;����l��Ւ_ѥMf��B������F�I"��7mOA�d�\5'��Q4i�l������UT� �%lmA�v��|\Ԩt�A(�:캿��s���:#�����/c��T(;o���4�*p} �B����<�9��j�%?��Kܿ�S`�C�K9m����������{�z�|?��|xƯ2����8��Ay�=
�ߞĚ��_֎������ǲ��]Y�x�6���V��T`���W|����xmPv���R� Jd��/�V��4V�-V�\$�qb����]��#�c���*dU꬧ '�K`������u]%^�(��>N�u2��Y��v�P1�}�m	տ(mi��jBH��( �O���n�n`��� �p�$�g�Kɫn	\��E���{^�������@��љ�bF��u��#�����]\�q ''��f6(��i�}��EM��kG��)���	�����)͒���,���ߋ}����Ϭ��t��	S�!oJլdYdQN0S�O��|d'A��jٴtHc���{����'�
0wwt�e��(� -��6���j��1$!��Ap;Ҫ��5H�<��4��A�^po ƑO�e����	R:5 R{:A��v��8�)?���^�+���a���|_���f�؉�;h�O���>�\�X���3���/o/B�[`Q}�σj�����[g���S@�̽����Y
y�7�o�E d��@[����5��jf��O����}oU��U,B���G8 ��ܟɫ��$��`�HQ�|wYa�lEPl|h���?���&T�����Q�N
<�.v����%��tf�ٖ����E.N�`��ǈ"%������CEqD(�TD'V*k���]'���n����n�󺂢�%�v�2�n�aM�D����
P��jmg���k�q%��1�#��`�M����L&bʶ��	�J�,��V�B��� �r��������$	�r{�Y@���:��'��&W�6��L�~_Q͆��Q� ��oܷ��Y�7���7�J!�޹�� ����6l\GU��������d��_3K*2(,��ީI&��)I��M��gfg�I~*���{�Q�˹)�s�:"������T���u"kDΟS3��ȗ̮'|qu�'U)�`!�jDa�q���B��c�Q8)y�
��\��pq�+M)ϡ��֞�o��_	����<u�����~��t��%hZ�����;6i_�eq�6�Z��VW��⸺_�����$��7Y��|����M�Բ�3��ހx�ڤ]����rV���/�8-Fgfdd��. W"�/��GV'�걆cbO?-���zdr�p*Mfeff����1&%f�?	4x����O���nU~��}{�Pb���Q�_`�G�l�x�,��IĽ��NZ]N�⧭1v[��D���v����������_�l�À-6�m��nx?�O1Q�)i�:����W�W�{S�/jl����a��h�6�(�V�;cAk9�l!�����|H�x�|���%��fP�<FtN�#V����5`� ��g�çP'fF�*�����|��v�#��KY�������uP��Q�v*#�𩰜������*tB�!�"x~�/�W>��'y�n<l�x����Kw!1��|���ݼ�l���~��4	��=g��	�5�.�j�����/�W#�K�}u�p�:�1�5�;0Ya}}�ZϾ��s�H�s|5�B�rz�k|x�nq��K"w��xBrk����ҳp��H�K���E�s�th	�����W��K�	8�#Ww��.g�Do��]�l�3��F�S3��_�H	��NW��!�7����#B� �~VUM��)E>��C�|U��A�����&���"��#�d�kŵe؆�y*���Pc4$�4��A��w,�̓���*��7w�\�#��el#5�V�����d��e덓4�ſ��Q�Y��6���������v Ų��Z��K9��YXe��tʊFJ�y�5�};�y������V�[X�A�3�T-������»��Xo��DC@@���%���fMS��{;OwK�v�*|���������DœLyV�ݣ���(��JuO)�q��O�<���\ZX��!&$Ԓg�}O�3R���wn&��Lo��Jz��歃������q�7`�P�� q��q��Һ�1Ew 2>m���%��'eT�հ"�@T�ЁTY&��	�1�H������ӗY�iU��6I���(Αc|�Cr�nk�R4JU�"�����6��(�+|v��QewQf�V�����%�\­�s�Q�-�ʪ�����8x���i�ŗ�� �B���;����l&a���6�x�Wg\Q�����}檥��v+_���4���z�x���xjx��yJ�R��V/�HȶK'�b0(b��全������QO_(2$���Q|�ۆ�a�w܈���J��n��}L��E_|�sń�4U�o$���h���x���J�5�1r���o�.v�OUe.��؈y:�qC�u��v�v]t���iz�ųq�/gB{�$PIE���T�6��o��(D~,�kg�� �&8���9�� �e0/F�	#��>1��=,��|G��w:vKH]���߭���s�^��G�M��f<�XH�$cI�'��dz�ʯm!#�88��z �䌬�����e@�!�o�x�_��z�^/-RPVۇ>��6˵����7�4b��!�#��+q9�!��i�Z�ܣi!bꙮ��2�9~B"B���9T��O�|M�xӮ�^� �k��Ol�#��)D�`�a'����PJR�92ҴCC��DC̸}�W�����e 	�6�Gr[�y�<���k�9��q�e#;��I�X결h�Uٓ�53�O���T�`��J����Vd^�����{�7V�:��y�,�N00d�J�Qru�>r���9��o�c��m<(ι���G���|�C"?�������k�N�φ�M�i�[=�(��[Ea�u�����m��9mV�,y|�^��0_BX�B�]YC�-�B�������w+�i��9��M�������-Dw��+`�\\pn���N�!�x�#��bznz?�FpD��U�ehu�,����z��ϭ�:BxzV~���?��rf\F�LnG�^lLLiz�w�����WCLa����\`���+*�%#��W�.w��ٸҤ0���������IÛ	���}ec#;=�7�6���xS.MY�w�J8$��?V0$ b�G�\D6���TJ%mR��GK��yۃ�L%�Q�Ԋٺ��?�*�A��-W��:��L!��pa9a�l֚�f�P���yVh!g������705��
�J�#������J�n���D�N
ulS���qO)! �|J#LH�B�;7�2�Az!*��d\g��C }�R�ӥ�[;�(�9�����pl���1!���s����5�fY���lk����&/�Z��x��!��_1@t�&��kd�q�sv��{��>��1���P��(Q�2�JOP�Y�#ӛbd�98�)q���T��l	�L)@ZY`V��sV@�r�ݦb*��Ӥ�ۼ�~�t�nWEg^���F����&�ĝf�����&^��k�r��й�'�ז��m'���E6��n��EE_q����ϟ?��@`����|�:��y��@��d�:���Z=\-�V���呣^�H/��U�-R�]�6�$2�zEp�R��[�l�[j���n��$�dx�%#���g�4,�Cxqvo��m�������5"����C�=�B,xR�Y<2R�
	,2�2>�Gj�+��z�aq�a��%{�����:��A�X���ub5��l:Uun�!*�9�;���3]�|ɣ�뾂�Ѿ�z�U;�}ٯ_��v�	���nk�ݕ����kʸNu�	��J���O�CBoW))X��y���h-�?�3^��Dx��W �4帒�'y;5L�''��Ԧ���5�Þ�k}�' ��P�z� ��(�$w
f��K#�	��`�eok 7�^�ps(V^e���s8��E���P␔�=��<�7kMcljw�-?����h""	�6�s���+��GH�'ڣ7s�{ZsW���A�)�i�E"1�9�ʁ��413ӆ�}p��a�%=ZkN(ҁ֟ª"6O�n��Wy���9%�|MMC�U��Q��h��C��D�bl�;��=�neeR��ti%O^X�t@�s���()�/�3��V�A5%/]�G���2��ssܫ��*Z��a�:���Ok-N�xg�������v
��.,�[7� I��ݾ��z�3�v�K�����ua��-E����Y�YvKt4�Ȑ�=��_(&�Ot�g-�h�,�.��Z�Y����+�����5ʊ�WA#
+
��C���^��Cm�[+�U�_[Ń*T�:��S�~��U߯_���4�w*!�IE@iY��EF~Όfܥ��J�,��89�%��Kg1>�5�7��
cn�</��&I�uot���������F�ɀ�T:(��.�&�UE��M���S�d��(�6��,�7똋�?r��ai�c"�H��<�����-#������#�ړ쬠���A
� ������ �]�ugO\�"���2�@5E&0d��u����dR�6��g1[
d�8�ߣ�r�)˲�t�����1�$��J��9�MM}�͹���鍅��������9�ͩ��]��B�o����c�@�����4�H�er��mD)���*�M�e�&U2���z�}��|��6�w����HM���C���)�l~/����	7� ��*g��X�MS�C1�����C�|n�Z���s���-5�$�HA}iG���[�5�c{
��(��M���no7\W�^W=_6�b����b���Bn�y�����d��;*O���me	ff�9�HJ�Ǉ/����!S6fv[h�`��'�x�s���R���o�Uo�5�1.8f�I�?q}M^��u����B�!�j�p#��14N[���U����Tf�����ɹs�����e	$��ښuF������_�ؖ5n�{��$�H!z_k�aH\�� ��Q;'^�������p��¯G�}>J�A��,Dq�B�$��p/�T�7^..��1�H��J��J85ʄ�r��<�:s<|�+�������veFH�I{7�.�'�������-�������t���_��r�5�1�1C$��n���
�7ݳ�P��_�%*���-XRwM7X>U�)Y�?���`��tVD�-H�Pr�a�EpL�����c[�O֮�s�2��k�Y�K�䣦;:Q���(o*��c��,��=�N����e=<='8o,l�s�����)���6��6C�W�@X?AX�<�N=ApX9k�|&�+ۖ�#?G\�� Q��boJ�6S��+��i�%000��Z H��JɊ�=��RF�.�jV-���qzm�d�,�0[Y?�z@�H�R ��}�������:�X�t������2���!hOU�f�
�S�
�'�&�6�:
=3����%�~γ�0B���8�, ����$Ďx���{*k@W�n��� J�����̝7��2KkH�
b�b	x��!~@�����x�9��|a��6�&B��dv����娔(���4�Kǉ��h���pRQ�c������e3��٢�D��om0��F���A�����r:��i׉9(�fT�?�D� ^^�ӷ���F����r`��������d�BX��;(Q�!}����t/+b�O֤?ӶAK�rt�e���>1�Q����++W;iz�h�^+�NFX�4��Т�7��c��]3�[�+�By�PO	5:��8�F,ʿ�٢	�m��}&�Bpg�	mk{e�\�;����QZ�$9��bW���	�{�H!��Z���Mф��j�ѡ?�y�Ie��Mv��3,=27̴���6 �[<4~sc��F)]gX�[���ƶ�8�d7|�3�.1��r{pؔ�بD���ђ97�F�������8�o� q���2�Rr�O�2�̲�D]?�9��Q����o�����5���V���#%~�bT�=0K�x���2���(S����G��w����
-�i����^���9���n���o��}��;+�n�R��Eϙ�y��R�*��oh}�v�dt�f�e��{�լ`٩ �us�E��fgm�@Q�r����"ώ���jeE�da���y�����:���3���%N�7%��'v��f�;$���W��0fW��)M��0-E�{��]9�iHK���f�إE���T��sK�p]���A�G�#6����:.�����f	�[=RS���-�T@�V��Vf�vԃ�B
�bE_2�-Ə.+��E�i&^6I��5��(��28%?��IaKOi�`���_,�뾅����v��LF\��8p�S��p�&J<�l�YȁG�-��<���8��%�����#���+���ξ�y��8.���R��56\Y.,D����C,�	�:�T��K�v��4B~Y�xn::9�jN�,g����Sm%bX^"q���߀!,\\�g�������Xqa��~�ك#��|A����s:�׸7u8�s66��R�-�����!::(YHK2�[����<?�(����O�֙̉T*~q�6V#����� q��Ͳ�����,��$�^����P�:6�R�����fR��7��rmWm��݁�<||#�=�<-���1�7,��K��9�>k?G"���
���N���\��a��j�-���%,r݁��뻓E��@b��h������n�E����f�E�5H2X^������r3N���l��i�88�����Z��}:o��{d�ǘ�v T�|E���������w��/O僌���G}�\N#?���%C:�lG��`8+�}��'�~����mL؁cݤ��������T�v�|�T�:7���DQPbH����DZ��(���|��ɏ̰�J_���Aʞ����~an��n"�h״yU׉v��dO�� r�4�h۩�d�ԙ+η�n;����V��C�!T�6g��YًZv�������4��~���8ߦ��׊(
��R�1F�:�kA�;�!��f]����4�:�6	��ş��z~D�y�v��t$5�TB����NϷ���FZ����^n��=i�;<V\?ɸ�{���.�Y<���P�8��&�������K@��*"B�h&_U�����v� ]���y�L���|�O���{x������G��kjLF#~��	��3c�ss333CW��={��s/_�6:2:
|�����(��������S�Ν;;rmxfz6�����R��T���ݷwo��5fk�%,lY{7:����]�Ov���dl�z8�Y����F�V�����V�%�k�T|�@� U��k��]kD��55��d217;3>6
�6��h����P"�� S��KPY4����8L��;'�˦��j�j
ǎ;~��z�N\ce��d� �rk�`0��ew��LT��f}��Tj)�Iga��.2ŕ�W�]ay�kyT�U}  ��?C�ݥh��� Mֻ�ʿ�*�7��ʰ�l�����1�:$5PTCCC`�J�]�'�8��v��'>18؏@�F�1Z}P�f[�D%�@ߛz��Չ2���m��4�Wð���)ډ&�'?�I�-M�< ��$��h�����]����1�:W���z㮚���9lo��j���t~����;>K�B1�u/�~�~>�js��{��3 w���2�
�{��1�y�[��a�<���]ݴ_�q�j����N���|��f� �����Q�Dk�7�Ƴ � Qy��۷�nvj���{%�R��BUCє�H����sO���ߟ:u
8�7�x�&P��s}���0�`q�v�m���*��Ղ������}6��=2���JMMMyJ�l	��1r��X)�>�8�����W�^6I$�&�\��-a�4�Qm(��>2:-��}���<ߴiP�G>�a��;���`o���n*\����C.Q`Np�	��K���4���K���|���*;;�?%p�Պ�X")q�*���5#��+�3�xlff�[*���8&�5�1Y�v�ޅ������y+��ؐQ�-��Ԯd�}tq�9B9&�!㯫��%'O��x��O�*4��M��T����}��r�aV��*�j�P���/��<�$$I������P�2�i����� ��'x
2����܊�-A����b<�֬Y�����Y�v�uU]�}�͆L#_�F�(��~�3���V9uܚ�������.��&�GЭ8�w�F�S�p�=�*MD���P���P���뒉��z,#4���@�� FZ��k:�����AKB��6>��DCA������"����������شiÖ͛wl۾~���������M�LW���b(A���Vý�5B,[*ۄ�􁜛��es��}wm]�O�z����կ*v\q�m2�38�"�s������~�7��o}��سwwggkMM4����H�Tȧөً.YZJONL�MO�e`Y:�hT*���Z[���uu�X�: ȉ��ɛo�55=�355�ZH�2�Xj�oرs�}ǎuvt`�/]������6�]1�̾��Gd7���2�[C�zJ��J&n�hJ@|$��I�F�ڵ��뿾{׮t:�P4��qɴ�b����i�D�"������D�����k�pGjZ (��d����!��P��ݸ۱c�x�@%��
.\LI�&�0�1�=�ɍ��,T%t`�������NCX����F�����[xW#���v8"��m�l���O
7��4�ހ��]�t7��v_c��4E��
}��b��b>���x�b%xkt����n��k?�яA��e��<����qM�P m[ ��ѭFr����ٳgΜ��i�������z��G�3����_n�($)W���L��q�a�P���L��>Ӯ4�T���;r��zؽ�R`�g)�q%pP��g���g��ys�l�S�@N  m�v�{�h�1�ƍ�x�	�㜺̹7�5 _�����C
�}�A��@��~�m�A<��n Zp��?|��Q #ud��@.�!B�	�jф0[)¡�A���!�]WW�ɓ'aQ4Nq���j��&g``�Oԭ�M.�r��fٻv0[��ٱ�E&i�A���O����'�5��0�{��СC �j���7�7]�c��0���+^�690K`^<�^�xL0��Vj ���n��8��=�{nO'������H�y�)��/��28���م����1�i�F`_�D�F�y:N�-��7�����@ɘ��Ǐ����].�((����ȑ�w���r <��4��L��F6������{}�|9�����%;~�U	ޖʽ���)v�X c���� H6�ΊFb\DM٠�Ǉ��K�M�H��#ێH�|HX�l*�d�( �L�AN��LLL���}�JY��V\��
"Y����>ã1 g6���Ђ&c����h���t`7kB��j�N`�;�	L~��LNN*�ܠT�.���P����qڻ\#dw&���.NU�Z&Z�;,��jh�������ۿ�������ݼySWWg��C}�hM4�LMN_�����K/-���� F����\���ΤR���[��2 x����ή�u��uvt%��u��%��:Ss&'.��7�G�RaQ��R�p(����%n�ZL�-<��7�����~�[�R?\u!�"�r���$Mʢ���������������3%7��ј�TX��6>6v�3�u�ʥ�3g.L�NGcɆ���D}ך�۶�����������{{����������w����74A0]�t�����]�d���E0��;�����0zmxjb,�C��7l�9���>�_��k�z�N*�=9+I:2a���g�'�LG;�W���y=��5�Cw#�T�P�*�s�njUR\r�� ��}�/|���D�S����#�a���BB|O�����.@:��!���40e`41xLd� � �	�	���7��U�Ȳ���
oHu0d��6�Í�6}����Q�PZ�|�=�} ^�,���I����������J����s��T�l�yb#i���Hc�4;R�0<4�A{�l��/�<=3%�*M��+�b]�E�X��a��2��v�l�sdZ�]@��&Ʀ�f�� ��V������/[^@�"f/&i�bv�-9���K��49>K��Y4[����	�kj�~��������A�0hկ��ƀ��Ճ/hSqw&u���]Z��P�F'Z�ŉ�~��70͎�:K�΄��Ї>t��ac}ЗLM�_\�F�.��!k@A��8��h�`*�4a {�bbe"�Q�'N\�t�(	��j��ATn��G?��{�s7�t:f��~�i�c���@Zq�,�L�uT�"]A��LNw����W��X��_���fЌ�?�0130��?L�&'G:[�1	����N/a��B-YW�D�^�87I�E��9l?��+W�0��IY>k��jU�k��}��M�6yz<hS-�!���i{�Q�y(f�vGʨJ>iL�s7J��ٝ�(.m��W^�es{�/�i��;w�:v��;�<����*U[>{��d����/7%���q�:0��с�9a<���,�&]��`{�s�>��/(��7�<M~n ����>P�&K�X	k��G<�t$��4d:C�M�or{��#@ҩԢɊ��B�1�Ⱦ�{{�={����}�#�Mk{�� �c>5��3[���,�p�Xʘ��c�����^�u��a׍�I$Sׯ_�裏9r4��f�#��jv+����f�̌T��^�%���er�����̱
�����%fZ~��ߔ���k����9��Nҹ�:SCꄤ�A�Nq<iK��}�<���@�/��\P�*(����þ.�ll�����ԓ��)^CK�ϛw	Ah�6n�|����0 ����B��t�O�3�<��V3%YY�������OMOMr�HX���b�L[AS�'��MkX����������T%�܂��n^�jX��ή���εk{ggR��t�M����K�T,�(�qcv�5���u}�p=�S$-a͡��пz�<SSS�idj�#���bo[�W�����;��@��Еr�?��'B�q��C�á �l?�R�L��� /�ؾ��{�~���C�ֻN0�Ƀ��hO�7��9s�ʕ񉩅T
�&�����!MO/���@:�3�sS��S���B ����5�}����?����[b5QS����6�X�����z9_�2� �����:�TjæqV����<��O�F��b)6�e���H���c?��������g���L6�%�Tv>��x��;o�����֞Ɩ�޾���e���2e�`՛.>k$'��������'O�<}�4�5����B?mذxbvf
w�FB��[�u�޽�������_�Ǣ�Ppa~�g�nI9^	�W�M"<��b!��d���h�m��׮�.,�¡X����wPx�}M�	�j��=��-�6j1��K`6�&=��*��� ��W����655�����u����lO����}*�Pƶm۞�γ�H(D��rJ0���a�g��ͱhL�k5��Sts��ZXL��L���H
�lnaa.'�PIL?O����9M� ��EʇE�,�/0//�u��+Kٜﺶ�>^�K���1�YZbPvy�t���g�}�������v1E��0���hnn�I��W����K����K$�x��۷]9U��=���x���4>'��g�%scjj����t
��M0m�ɾI��?@�Lǹ��"J�r8p`�����ƨI �.�Ju,���Ơ���3i������T�]]k�jk��,f/Mb'&���d&����Q�0����k�a���ϔ�
`}��9+H��R�!�\�)v�'���� �`����A|�v����|Y,��C�`��LMk�MU���Ч���M�k��b5�����8���(�)_Q��� �P0�52���4��P��s��w�y�4�-%8~B����͛7r��:c��k�'R,���V����bz�d\�4.D�Ov^.��DdwZQ~�#��9f/~��9�b�Ӥ�i������\)mc�`�z�����!h��x���eIV'���{a�;v� �?{�,ۅi�lV~��.F���
w���vTQP�t+"�n�HE~�^,��`7�� ؀��Iq�(-sf��[�n߾�駿)�-=��>�>g,�Hks�[�1����g�Zhjj�1+�����V��4;۔�;8�l��,:H�300�Հ��J�&&�9��v�R1[��t�U�0�M��E�@}]=�%����BB3�V��}�$7JA�R�TF���R,inl�\����+a���
�
���T��&�&��	)hvy�h�������Jj��?h�-wZZZ!p����x'�Y*')��.{�߿��]�4��Cͽ�v���|�X?A=��Dm�	:K҂�{X�ش ʡ��Tq��q��*Ԙ8@2\7�KRtXv��� 77�;�h�y����+�-�ko�Jՠ[��J ,4�:����꺺q �](����L?��ʡ���}�Ɏ��Ղ���o���a�`������d��bjf�J0��l���W._��!����;�ȱ(�=q0�-�⃱:37;=� B
�xM�grb*V�hn�lk�O��|���5[�m�w��/}�K/��=�+��*!����T�K_9��#	>L��0q@��<��]w��6�n�� #�&3!��H4�����|�O�w�K�q�'"��I�] <s��##c�p��mMGGצ�ہ�ZZdWGȉb.c:�d�X5B/�����dC�tAO6��=x`�����׏_�p��嗿ύ�Qq��������?���������׋�)H������d�9�H�L�v�?w�����<xb�����g�}�{Ͻ04|��O��V���1C�?�ğ��"������ЧN؈K���Z�v��	,
Pī(�t*'X6o|�����؅�{3�o߁��VkKo�`�R^�m�q��=]�m�#I���%�`�S��5��S��u���ɤ'&�d��7�P@^Cm� ��ے�;�$��֭[��Ԥ��~!2�꒐|bKk���������M��=���M0HP�`W�!,���>;;�D�\�����x��[\�x��������U0�Ψ��0�@c�������f3��X)"��#�xZǟ��RCRrS���\��@u���+��/�ȏ/�i� ��5 7_����������L��wU�N�vf��ˊ���,�$^SĄ�EH�i#L��� |�Aa3^Z�þ�l:�-V�ȑ#���w`�x2�*���Y�n�@�|��rU7VKS
3��P�����������76$k����Cٯ&3	1���w�W�򕡡!헠�&�7�#����{J�� crb�ԩ�)fL�>��)����>Xpv%�K?p�K��̩S�t%;��b� 1�s51E����徐�`�e��T��6���bv+IRZ���@���C���z�9ooo��LmFb��ڨ��	��5��%����>��ّ�Eq����7o~�駙����4���M8��+9+yˠ���'1�Eh�T����LT~pbb���X`�,��v���T�~˖-���}���A�r[6�Y__�Ě{;��]t��0������0��,�f�l�
�T��N�׷7�b�o۶�P��T�'����&���78؏�`c�y�
xӂ"�B�$b�~��g��V�Y��Y�fM8$ilb8��Ǥ�a���i3pN���ebrv��q�NgiE��p�w�&�f�J��B���ކ�Fj�x`���|�;�^�ʑȹ��V���A��-M;vl۲e,g�jKZ�m ��y 8�0?O2pT�(������:Zk�%c�uL���;>ɶ qb	�R`ϡ�+��gz�f?F���V)Y#��4eBh:J�L��]ɀb�sp�L`�;�m'�}#Z�&��k]�y��7~�r��VЊ��2Ĭ � �u}]�+}y{��ٷo/4���J$�͝3���\�� ��l�gV�;�ɖ�u-�Ufz��a��2���B.�+��~�l����I�65�Fc�斆{�w����k_��O�u���X�1��W*��t��N%MN�p <9� t�O����`#}�f�<�ɏ~�W~�W�zs�L:��K�-�r��3gΝ9qnfz���m��]�m�]��_vzznd����|CC]WG'��B�T��ʽ�"a᜜�L�>�����#���w��������_����۷o?{&V������;���}ntl���!��P�ZDa3��!V��^.Z3B~��m�?�$ ������s���������U�;���C�]6un�
"d�C��΃�Ғ4�q��h��0�Cz�!�` ��Ov���355����KM�m�&� =�� �0;��^s`�>�ӽ:T�����S_�ȝ++��'�͠jV�@�www�`-���PN��$�LLMN�L�8g��ѣ�a.�8�ԡɌ*�^X>�bmosS���Ҁ	�b���x� S��+;~�0��'O��? �b�'|ǃh�{/��T�� �s�`���˨g9�a6�,���B�
��ׯhin�������=s|d;龾>��@�E�����)i=r� ���!(��b0��8��ŋ�#XЄ���t""��d��PǴ;��Ȍ��"�3䏄#XiV�B[�Q��di)e�x�K����2X�W^y����f�/z��a&���m��tw���#遛����n���d*.�5�)-�&&� #@�6�c)C'b���ӧ���c#�.P�� ��'n,�������Z�*��؇x��g�b���+q�%X�xq19��J�v�&�3=9y��E,:`d2�.S��5� #'�&>j������h#:�:	�#�����/c�٘[H+TΖў`s���6�e�C����.��a0~�;#�v�ҟ'�ZZ� ��A�ґܞ
��}X��!��13,�by��Y�3��[5�]
��ō�ߗ/_֍���1���m�m3@�)��V-��>�R,Ig���Qn>�s��Ij�''3�'|gG@��q!�C�WW��y.�ʊ�|�m���}��\"^��چ�Mۺ����-B!ΐ� ̒�I|�Yl醛���������b�*n�ƞ����=��!��=Ŋ�́{��%LB�5���/]��U����%3��q���,�A��b�\�y�H_��Q��.q;f������rXȚX���{:�ڵ^n�,��A���UPcn�L���aj����K�x⦍[�6�C�mWv �S��eNѴ6��9���������]G�/�K��OA�;�ť������q�����2�+݉�EcK�\��h��hhl�b���ҝ/ ƌ��;;۱CC�5�2K攊�WW�J��u���O6�in4���]*f1qaR����M}P9���s��3�a�&�!��6#1ُ%mޤ!�,S�����
���Ǌ��&�E�P���!������z�СC[�l��� `̘B�4�Z�zu���s�E������۰	��(u���J��c45/3�tZ�;�Nr�vm����cc�3X����ơ��8��斶d]c<V
��s�=}����k��:19Vt��p0oZ��n+9����C�|(��E�̾��܌Ŗ�Ko���$�ӓ��V����L:�������������>K�𚑠���&�F_���|*K��]�e[#�h�����&��{6VI��%�ii�8����Yɭ*}�+>&�W�Y��&�;O;�2���;�l�����������㗾t�̙�{��|���~f����7�����~�w&&����x��X���+ƣ�Tzq����y�3��-g���dT;>��Bjǳ�r�������wo߶�oΗ��&���z7(��I�BF�����"s������̲�"��#��z/�Q܅F�[�":� �)|35>q)q�����Z̪��q�ȇ�L���vxcvaqvn!�d�W�c�1OX]]� xL�jr�`0�zP��7o�0�NE�VV��X���K�)dǉ�zz��v���d��	$�EB�
**��C�����uG��Ë���&Xڥb>��h���5rm�����Rd��ںi�f:�g�d�H�h$RW[�K�fg� }F����D�����:�Z��-m��P1'���P���p) �#Eh��bbξP0���8�c�"QQN������~�ĉ�8�k��X�� ����ݯ���D����sܴ^�+4�D�z��lݴ~]_���)�K�} s��L�P�v��j?o����c�=��1I0��������o�v❷��d�ϐ$��um��2!���dM���ulb
�tb��)��+Y��+�M��(����曰_x�\q����p9�h3$��GF_����ƵP6 u�Q;yX�=�����`_(�dM��@��' m�M�yV4b��3cA!?Fzƒ�n׬�Js<c���� _�tujrk��j�o��/����K�=��Ҵa���ߒ<+����A֨����YS,0P&f�!�D�u���ϝy��7�:�w�ŵ�b[����`HN_XZ�$$��N���4E:�F`�,U�!���J%�Z�i6�\6C<�CRW3r�Xx��Up�ƍ[�fJ�{�J+#�0�ݺm�˂�M����d
�j*�7�۴��Ņ�X�P����']�r��A<1����D�|����4�1�f:���QQ4`7��
�A�Ν���'Vz���>�Tpa�6���x@J��D蛔z���	,n���0�|��D�&4љ3�����A��6Ic��3�B2Ƀ�a�F��ա��kx2����������߀��l0���}eb�� 炴 ��J�B0̝�ˑ7zEK� �Ϟ9�j�B�! �:�4�?_��"Q���_�����^]S#�1����1l�؁9WL�]n�Ln޸$*��x���<F�@o������cx��1����k(,�,xp)�a��z�!G�7��	���q�n1_������nok�?���'�O@H|[E�R7�/udd����,��$��q�~���>��[��t����\C�LxVB^rO1Hڼ�AQv�R�%(hkl�r&�����ΐ�E���u�	�����j���!�AK�bZԘF<4��a�Q�X�S�K��@�b�8?�h�-�y����{�9������>*�؁��;�c�.�"�
b���y�)�W(mݺu����ݶ�t�,1
SN܍��&-��wM�V_8GE�6�6�6u��p���g'�F��gF�&'�&kk��}P�M�m͍u�۶�t��6�~�+_���}���%�n(�\�����,�4(�f_J(�S�_PP\�p�ʕ+?�Ѝ�R�Rް��ʤ3�6������/��/GbqY�B��]�8������7_���w�ڼx�7�L����L�)r����v0��	&�� �%�&�
Ģ��Jame6��i�3�O:|������Ɏ���g-f6�J}�������ۉ3��3/%�ъ�"����w���9��u5J�-e|咰���@t0 ��e�)O�K����E�(P��z
*l�Ȋ6һ,��I7��F��a$H>t6�è�����Bj��k��A�Y��"bQ�"��e3�0te��X��s��*��K2��r��h�l�%}H��n#0D��B��`~(-��M�(@f��٩��.�Y��&ZGp+��}����<��891	K�}���';;;1��IIWÛVoQ����_2��~D��+���.wQ0M]��2/��:�l
����z������Bj�q``]}}^�5�H��� ��6JD#����|tN�f����NMB+,l����J�ϩS�~��0�
��F>?�(nȉ	�N~@�~������u����S�)M��*$%"3v�����y�׵#���冝����H&a�ry����[�`�`r��Kߤ�I�qCi�]������ ��_~����c�AV���R$*���+��\cC���4[�\	�F<�e�a�E�Tj�҅gO��Eq��Y ������nI8�׮MNL0�<2 p5���Μ9#ӤV2�������Ż�?��.���K*�X4�YcV��z:�h)/y��L� ��J�4��ݽ�8���N�=jzf�g�qx/���)��#Ѩk:m���Ў ?L;wyT�Tjϒ���ֶ��eOOe͒�~�4'O��m�FF@*�Xxs+�o8kvv9=5}��񎎶�{v�`\Ǔ��߿s��7�x��p0d�\+�}�j�%|�4Y�2P���$$��90�|���M� 0K�)�쨉�C��ʯ��V�x)<T|����_���ȖĲ�����{@�u�g��^��:�n4B#�(R$%�%��D˖%���x<g��{����9��Y��0����3�ǲ�$�E� &� ����Xݕ������~h&%Js�UwW�w߽������grA��!�V=L����`+�����B40��5H�fzx�r�N�:��MV�u�^�4;����F�QH�,e�Tl��E��`Fɖ�ِ�v�kڼ4ˍM<�	����e����F��z{k���˗''� �d�I����*�fZ�0�@�`�$�^���j�dӎ��D��l["�T�Wc�R+���j�T�*`���2��O�4y1 ��6��[/�����@�I&]A^�_'�c1�P�8�g�a�]��<��E~��n�p��:�����J��+�DT�]���I}��'�	�O}�ҥ7.���Ɇ���tZD���	w�X�Xʉ����5�1��N�ۓ	RP�b@�6r¦����>
�b}zj���ۅ]C������}}�x�ɩ�����TY�l���}wA�R[X�x"��:��e��vl���a(�a� L����l?��D!�W^/���|��%,%�sX��E4O��6��N�>�������g1����?��4���*E�W���<66�g�޻?�	X��8���r'O���so_��=�ٕn�d\ĕ�LO�ېգ�q�끛M��e�U����o�1����(��^-�� ��\Z�<>�k����p��7��������Ï>ry���X���.pW90�is�@%�?��a^Ӄ����?&)6��y�PC0�����P�Ѭ�5Q7
K�q��so�y!�=z�7�ٳ��=I�D��Zn�b���	Z}T��> �j@�{h
�]�y�(�`��m�el���������~��я,528<q�L4��wHο�����Ξ� Z���֙J�}-�·<��N��rgcĦ�;�b��O��4}��$Lq�?�
G"��Pk�T��|�6�����~:�9�@�I��� ���$��ȗ c���=K��J�|6*l`6�iddS�����6���Ū�J�S��z�4e����^1�ŽtÒ(�����j3ukyqivz&�j�'c�E���k�&'�@5@S���`κ������.B�TJ i6�|���O¬��䃘;3�ZA-�C��U� S�h-�h����Y�~�tj�"�?@���ָ�abbbxd8 ��i�����W�-�Q���F�dr��H�c#�t�E���dŒ��E�;�5�Ҁ�.�r�����,> ��NwD"�"�י3g���(�(r0�����d ��R�*�;Н0���nz��������En�����brp#A9t\��"��j@3 �0����2p�M��x�2���9p����Bw�qQ�	k��ȴ �դ��r�0��X������ԩf�&���PΜ]
1CwQ/��l҄ޯ�+�Z���x!u�Ƥyf�h%ߐ�$��nZ,���V�N������ѥ���a���0 \��mE�N4c[`��˴���S���$��q��_���p6��5����0G}'�V���(C�6 dġ��<+a��azU�x��`� 1u�R%�������"��W8��'��d6��x||em����	�΀J���ͬ Pb�����T�6�_q|���x5'8a��.k-����MV�8}4?�L�0)c�w�>���axͦ��X8��SI�)�c:d�QD@ͱ2Tr|�����ʛ'N-�,a�b����0%P�|ɤ���).&Ը����\ƎhT��W��]�-"�0��0kv��1��#)TvK�'��M�"G��24i��F@�4	� V&gxxHqQ%@r"��RiQZp���o�aAH8�B�9��RT�E�,v�
H��ĮA*@5��+�����g����X5�*;G::�E�T�C�}F�@ ��X�R�d��Ֆ6k�z8b*.����i~|",�I��rpl���k�V�W W�u���^�����T7��<$�ec�H2W$_�V���*o�*��mE�l�"��#�/1�%��P�-k�\+���NYjոJ���Z1�"6�7��gϝ>}�R*�(n۶�\���`XWu�UP��PԴ���3�R���a{{{p=L[�8f�L�u6y�n��ݮR��L�.-�`Z��+��R_�Y��JJ�Y��9~) +-
3K�u�\ƼA`�(�/zF���G	��1N`�M/�mL�S�|�����eC��ԕ]q=�8�*��D���M��ۇn���z�b
pwb�<�e����\s �P,���*�����*v8��^�:1���r�3�S�p,.ZVQ�������}|�V|��7^���+6�eN������vfײ�=��~�a�O<����F��W%QG)�x����&�ʢ���vc�� î?u��OE��?" +
�?�����~��;��x�n6p*,/��Nͬ�?�ѡ�mcC=�t�p*��`A�DbQ��߄�۲[�7-��R�|�0���z�J�tM��n{�(������o�Ϳ����_����f��s����M������/~�X�2[(�A}-t�xo�z�ۨf<5ʡ�V�O��/�|��G����PN�O蜙�����sףG�BR�SD����(q9ְ�RJ���%���P�v�R��D A �b&�m8� \|���F��(r ��V-�l;���JU�CT�`R��i:tSw$�qr :���`-`����@���d���F�R�U��ٙ�����+�+8�n�P�s7��E"�յ�t�ψ�W2d���f���� �(]��%��ej_�X�cT���#c|<����8m�� %�� Rf,���.^łc�p\;$�&䷆�9-��ֽ4-A�-���e�q�RY�S�4��<~�����Ϟ=��;w477W+W�(i�K�A��j��'kX��;�p����oML��%ܫk|5  T�ި51TEu>v+��r� !X\ǖw�3�R�0�B���"�θSR@�[+-�}}=�C��=�1�1n���3D�}&��0Sp.��t��!�m��|�$�� ����/^�p!	1]�c�@rb�+X.DJU%ƓԐ� �z�&x�b���T`M��zi��m�ن]��Es�5�m���;���4a�&Ri�0V,�)��֛F�R[Y[e� H#��L�t�i2�NC	c�=����%�E-��O�+>��XN�M��Z%���+�,SqG&��a��K��v ���aTJU��4���n՛M�sr���&(y�)���h�L� �
q��*��u�@*����z�Ň)	>Ĭ�as���Gq��HP>8)��}5�������K�;��r�ׁЭu`�d*!����6�&�:55�'J�4��Y���*�sR�Z���H �T��e�1x��0A�G��S�6?g#S�0���RrL�t<	��
؞����?Y�)&''9"���U���NTi�h�^�b��2����"e̎a�܋&��a�kj�!�iC��j�u�?�|;]��x���(@I}������,��¼�m����x�i:L�Q��"#�c`E"1���aȊ��lc�e�	U	�"����;oK��7.>11A�p��CQ��Lf�ҴkR�&Ǝy�d3�l��0ވ��8VC<4¥M�yѣ�'�N-��/_�-���4efp fպX
lN��'N��xq
h*�����z ��}<���jH�em5��U������������ΥI	�"*8��p�6����TH�c�S�0�y_�{fcH�>'�*D`�@+�/&B��(���.j��(�ݱ����W�+���G������q�_ou�b�|�ԣ�p2h����?��[�-��,/�Z�˯���ݲe�]wݵo�>(9*�"~]F~]T|��vl����`_6w{.b"P�]������H<�ޙ���qV�Q�B,���+�5���z���+~%��۶�X)�w����x�_[�������B�h~*n����T�!7P��l���W��D�D�;��m��ʚ�6IQ����{�{,�}���6k�����g�}���e)��<>�3ܞn7�F!�'��"���_�r�?�{�c@y�R�w-&S��#b�. �(-��� ��-[�������o������w��[?<3���٥�?���l��?��J�	�jz3��e���l%Mn0Q��c+�Fu]�/�7�&͞#��0�D�J�<(���:p5�����ᩃ����S�n��8�ʑW\I�l�V����IGz�o���X�1H?��?ug��1�!J꯽�#Of(Z⚂NQ�w�y�믿>33��,�wuU�}�U|8 ЏS�G$2�\����ڵkW��%�9��|ɯ@�0��F�j�����7��ϰ�P$�N���%ѭ¤֨�MD4���}}CP�s�s�@�T(X��0�0�+W��tdH����` �C�ē1�/��=5�1�����()��T��E1����VȮ������B�O�i!��d�� q�J�RQԷ�������*py~-K$T0�l(j��1�ɑ^��J�$�tr/����]�ԳkyAD�_
�b,՛u�R�Ct�	�pE��p�� ִ��;�IM90!��H@�t�G*拥J�
,��������ކ*����h��o�*��t��Ck+`}�ږm[�����d2����'p�m5�&1@�#a��
 ��r܍�{�pK�B��w�g
��Lֵ1�������������s�@x�Jյ�|6k4W.oݼ����Y/�?;������܉�|��ת�2�Dm)+����E����X,kTPo`��T���v�0��63	S��� �c��u������` K>��w���B��Y�����A|�  L@��O�L�^�a��ǋ/2e�`�KA',/-@`ڻmm!�_�����"&Y!?�
Xfei	�E�,\�c#�D�5�gfqM�Ҁ�lVq?4j�^)�`�dr�j��k6��D,b�b��Ń�?��B)�� 6�;S]����rڶ�A�^�����&�<Mi<�)���E��ϫ�:.���=����lf����?��O`���"�a4cWl}���NOR�'�f�NO��l1���������>s� �����A�ـLj�Z�V�,��)�	��*���Vs񸾺��;��������1��������HD��YZ�+���0�:/nʪ��11X��V�)�8�DxI��[=j�XS�����lM�: ��^�;?5Q��Hq-�a�{��ʕF���2e')�8	u�k�E^h^_��s�G䇰O�w���cfnn^SZ������v��sٌ�n�\��U.\-�A�����/�cWw���k��e�4FFF"�0��JİS��k>{��H8��׉�*5���j��*;}h>�E�W����k5�f�o�{�.���H��m����[^���w����P!#�9��<5rQ"�e�����)]�k���Z�\o�5r��.�p3O3L��[�o͕a���֠���)�~hY�Ui)�˯�O.��d2�۶m�¹r�6x�R�����k�*�nN-�-"q��b�c�^L@�'�(�%�"�Nb�Mŧ�~���t�teu9�hO��`Q��q�4�[8>��f��\_�՛����,U���� ���/�Z@�Wj��P6۷����K08:RmMC?}����|�x�#�BS7��)�1�]��%7�	����s�G��\���*6�����-�H���u"F���4<��g/�^j��o��c�fgg�J'n�B���p��_��C����
ٵtǲ���$�9�y�}��+��v� �mK5!ڲ�>�s��zk_� �{$��V_X*!Σ���"/ΟH\e���Ǝ�KK+0�3�+k���D4�N�C!�5����w|��k���z!���}�z��#��60\KI��@��F����7�Y���d��p$;��`�U��[��7MC�bo����4�s{f�x�����y��S�����Ͷ�x�R���,2���Ź�Xg�?	�����K=흩d��� D N�l̟�a��^�f�a�������_��_��������W��{�����Z ���/dI�����f#�H�Y����ખZ��m��k�J<y>E1LC�4���Q�j�H�8��^?r���#G�~9�ݢ�j�$p�;\%���9�X��v�k���Z@hF�`p��R��9]8`��!��/|�3��VŹ��d��W�p�6���8�ax0�s�e�eY�E�0	,������ܖ�X�!2F��d��z�hJ��j+8D�~mymaa�Z��r�Ќ� ���yΆ"�d�R����2�Ç���i�_�,8�˯�1��!�����&B.�V:8��\��7��T�P(�g
��8����0v��_���-�2� y�M]1[�4\6qz�נ��Ү�<�9x�n�k��Q�\Mo�����"�SA��!)h0��gv��q��)\�80<��R�8��lKc�q���<.�r8��Iom��	HA�T�VƯ*z�Z�U������.G����sW.s�-,�s��l۶�ȑ� �n��f�������V���-��1 Yⴐ6�;n����cF#|��z��T��GXYYZ^�`u��7��M�==�r���-�/ �s	���3g�E�>Ğ-�L� �їq�7;;���,N��1��N\��+�q)@�#�op#H��-D�'ߛo���| ���~�F&2�籬L"")$6XY����i�,{>٫aFQ�L��G����-(#���@J��Ȧ�}AJ)�c-�X�%��J���������'�b$"�'����M�b�d���"�>NO�p�	?~��H��V�ˡ�9Y,YUhr6s tw�cj8n��}T���`ċ�o \��%��1�Zä���E������؜��.�Tk̩-)*�ab �\2�%�W ���`��.�1�����wjj
_Ĩ�s�����utw�֛TB~0$I���Dg��p+�C�\�N�b˳9�fr�����<�Þ��1*֨�7<������#9a���y�ַHt��h[��n��@t�Vn���tj ��߳gOONNr��$��;t�W�(��yG�WH2�	�_<$�J��	
62-��23��y�xY���{�ɥ������?��3-�3�t��])Vp���~fu"	��Sk:���19��¤�܃ezz��� ����#� ���64��	R�ʂI�}Ld���/HM�:Ҋ9w9��yDqk���L�!����(ˋ�u|2KxոK���T~�Z��IcI�b/CF~1�ȰlS\�I����ě,�lE�^�B|gC���� f˖-�|;�M�g"�fq9a�3k�Ui��OG���yJ5��-K��7 %�ٱp�#�*s��_���o��w(�{j
�{f��m�0�7o����F,�����	7~a��c�2A�JR�m�J��Ń�^{MW{���M�>�Y*o�t�ĉ`���ZN�0��n��Zn����\�e%˥`�h���=����J|m4 B��h�}3��s�'��W'���$�����ڵEoX�,�5�6��/���GNM��ط�������Tlr�t.����K%���iP�5�S���}dy�b��l�������_�g�y��۷���ٙ�����{�/�t��Ǟэyg�j�ƹ�� ��B�13!8à�4ѐ[T 4q��[�(F���x�h��9VCP�Ɛ�-�����$�m|)�n��8�{:��������ؑ[R2��0:q��8�z�oڄӁM�!���lf�4:�_dKH�jXN]!GE�UaI�a۳	��p-���#���
S�K���ܰ�
�������[�PO$�=���+*�X�o�����V�,%��/*�%X���6�ANQ�g�F��]I>�/,���ٖõ@�����m4��>wԠ�
mc�Ҁ#��S�r�KĒՀ�죬|G��;�6F�"𥉉�����D�.L%$F��L;Q͏�3��^�j��� J5@����T��L����t�H�^S�9��.㒷��\�υ��"%	e ��bWH���H>��� � ���.���{ixx�{�8��`R�~(�O�(����+hrQ����0Z�(!"��ǹ�PT�G�4��/��iӦ�|�3����!ęf�#��x��g�b0��GQ@���i66Y�9��Q�@���oN��S�q�ر���#�<#n�O�89`� �鈑P���
�]������*�L26�X�F���A�o,���a�a�.aB��3g)���+�I��#�� C��t�C:���#�{��0 N��]D1���B��*=!0�$��m����l3(����03@��!�6YP:���=�P�k����1e.fLN�T���f�x~�O�;��{���+�2�7��aQ�K688�[�9�8{�]-�������G&">� W�Oe��5`�4I�H�s{%\�Y�aH���oݺ�3�X�w����K/a� ��I�|},�$���)1�u7&i�b��'�8�YΦY-W�kT��9o�k�o�����c`�A��3�g<&
�%�������c��׳�D?"�;"y����5�2t��(�0v�U�Ӷ՛&��z��9���Vʬ���,1�����K#��W����ҚrS����K�/A�s�ݶY+��W(lT۴��g�|���=Ȏ'�m���,4�Z*��*`~�lC��J	����ǌ��d>���vu���2M�	��Ti�����0�a�$��J1LK�#YAq�.�c{�;�Z��l@�r�
� �vd��3�Lܥ�U�4�����山���tP?�&Џ��c���Qq��Z�Y�`߯��}��v�"�&����t�P޳g�}� 	�;���C@�����=1)eYg�\.E�c�6U	�"���[|�ocv�B&S
�aî@4i3L{td��;������Ǜ�2���U���+������5}?!������]w�%Ev�?����C��(܌�p����+_y��ŭ��r�ͷ���t��\�Zk��)*r^cM�j�߉��I���|\k�(�@0������?����O�����4nv��/������^�|:�*����5p�f#��{���N��t���7!��������N�j ?��_��w?�����V7�2͹���+�����}�m콋�~�!Γ��6��}�ʄ�B�1{#�����~�ט���m_�p��oQOk��JJ6���p��d��,X~�m�s�SV��B�l��)*7�إ�+��T�m��l6?3s�
��+��������8Fcrr�\����\�j��Aٴ~�շ a42��x��p��.$�g�nPC����K����Jh������(����.le�.,���ɑ���O��7j�X"��r�Y|	*ej7�DD�����D��w��3�qM�y�tL��1���s�=�� y��:�`B	<)֋/�y�GJ.��-b&�����Ć�OzK8�=�\d���ƬlQ �Ax��V��+����xf��;���Pa��=��c��>�1�KrRF�V%D��)�w��O�����G�{se��e0x_*����!�1�r���oߎ%&f�F���/B~X���zL�P8��()�1��lG���LQ0an�p@��$菳c��2�g!dO-���d��oq��8��ؗ��FG�a��kD]E�*7u���ֽ�$�9�KQ�t�h49�G���Z�)���,W�2NhX;ܤ����x�bx�w�f[����� f�Et�6�g�׼�>ǂ�'l%���Mѹ��p�á�����_�]ƶn�
�+�q;@@�3�iaTc`���^j���[�Npw~(/!��錘�]H#�3�衎��j�G^:̍\�U\�D�wvR�"c~ 0��ٳg�����G�{z���a&y7�)�"�O����H�@��89�)�����Ǜ�G�^<�5g�����>Zb��b�%9t�PGW',I�!�4�L�����#y�~E89��k�5�L�I�����a�3��}���`�B�+e��0Y 16��ܰ�D8	���Ŵ"�J���:�'H��VO-�j[=Uh}1P�'����ڻ�a4s�_c�l���g`� �1��RLU��������!wWݗ!s{J���ՑM�#a-(ܩ�藨�®k��������(�j���p�`�"�k9��΂������� �=;2D��c�RN�e��S�$Gb�Q�����rV���"��D�/C�≶�٩)l(�[ׄ�h�C%�u~���}F�d����n�?�?�`��W���B�$Â1,�џ��Ԍ�q�7������H�B��v��\�p��]������)H�	{��������f�9���ؾ�Dfe��%Ϟko��������V�z1s���  ��tc,������ӟ_Yοy��F�$=�%Z/j>�r��
��cC观,A8PO^Y�ך�d9w���}��9�E;?�Tkmy��ą�La|���?p��(�'Q/��.���A������g��`�w^�Ż���lPfE$��}����8y��{ �'�m ����ӿ������e����^p��U����`���?����j.t���#�~HS��^{������׿^̗��R�F'����;�V�K��Gߘ����6���82���9&�-qX�p.
>���B�8p ��xq�RhD�v,T9:�Aq���X �7(��X!���*y�D��J��k���LxV�:8دP]����TF����/����޽����������`A�7sy4g�ǡ4ni%K�NEF�R�L?N�j5á�)�A��J�墉Pf��^I>z�NLL<���'~��{ h<���2�).��6��.�U�Ȫ�En���YZ	i>��v"��$�<������\���<N;��`�egt���\`�i�j5��ە��� �7~�JeMs}�B��04�;�`)9�Ӣ�q����oA��+%�2@Nz�jӹ#��؅AB(���h����:uJ40!�n��xyY:�Om4LYrY 9���A�;�C�w	�ԫ�������j�9Q��#��-G��D���*�B���srX���#�(KzS@�nQ���&R�ȠvXL��dfp ,��9E�3�Dp�b5�OpqBr��[Y��o�Du����z��<��X��F�uWTN�Y�m�؃�P��
s���]�B4	2U<q���&!v�c���A6�X�b��6�4+�H��=k�gƬ���\�����E���0�<n��t�l^�<@�5&��|HѮ��lO������a� d�,^l^�2u�O8��|�F�LhO�Rׇ��Qd��`��"�D]�\��Y#�g�AʩG,���T��U��Q�YD�j;vP�N&2�hp6��O�ٙx#�Gh�M"3N3vE���5�X�;�r܌cnP�5��p �C]���b�ƾ������2g��`˶�W��2zc����҈�_�rLط"��ț�!�0<C��x�7�%&D���499�c޿?!GPl�5��	7�~�AI�'"�,�:��;��I�q�K��C��q �����+aqc!��V$Q9����tm޼:��ʓ/|���7�fb̺m֕��"+K��8�d���J�ZM`! �P�l�S��X>H��ݴiS"��驉]�)����-�<�����Z��iIա�����NG�9�Y�D[^�����b�@3c0*��"�c��Z|��j��}�z&���������8>�+L\�Ve�)���}�=��v�m�}������s&c��'?y�ؖ�P�����nco��#���f ��݋S`qz���3վ��T[*����7<����w�f�����?4�9��"IE����_0����^�:�,3��'λF��G����4����{��1<f��h���w�366DY�zUi�ie3k���w����n�|��>׬/�_iK�B��#S�G�oMh���}�V�?r|e�s���V*CC���{�P�tX7�ٺeT����z�����'�*�i��wcr�ך�d�s���/�z��[_?0`��o���ƍ&q�^��@WW��*_�җ��׌r��K�{��F}�㼿!`<�}�F3�Y\ ��s�K,�W���+_�
�n�9���k'��TN�j����6u*��:��Q�Q!b:i$6�DP�f��+���ii��ݎhs�E*�"'�qv,4���}���^��"E!4o6�����p���8�)��4j�
��˪_�x(<;#!�&��Z'>'��dG��={p)��z�qj�_|�ř��ݻw�c\ȎI`i�7��9��c�8!��	R,H�������a`c\D�,D��v�"t��١x𩩩�;���&=n0��l��z=r�ȇ?�a�@�o��&�+K��3��j
�ؚ�*(�LP�SƔ����&�1A�U'�p�cN��<�N:��E���\�sssO>�d&�<<<��qʞ9s�o?�g�us��WSA�0�%�9O���(���\��ɽ���d�����!7$�"�
1���?����_�����8����p���xv���ZA�[Ո�" ���9??��o4ukݷbʾV-�C�\5A,Nq|��7�خ�,<0\{��_[;}��ɓ'!�<�q�\\��p�n
�%�Ka	p;�fx.�i�Ø�gG�Y�P�*�,~O������������Z��Ҙ"�~�nL"����`����Ѱ��E��2�H��Ɣ"�@�4x��vw���q9��lerĀ3�8��_�ԧ>�u��q�cǎA� ^��叅��w�l��D�c��'�@�'�̘ ���P���`�q�	�?�;�,L�X�+~ɓ32:Z*��P
�y�����=D�3Q!B�z�F{��4Ƶ^�$�jkc�����>9a�Rݎeau����Q��Ik��Х���@	��\Y~UK���a,��%��XE5a���М�Alo-8l�W,;�s�����w�u��7z�g��гu3+��!�/����0�$�[9r�*�GL���#���y����+�S�Na�ש/b�5 ւ�u�p�5��a!��yn��0��<܂A�me{�&^r�e�l6��(1;#T�-�k��p,��ڕ+�|2,X[(6�$펮.
���K��N�>�^!��]O�ar�L�J �d
��4,<][[������9�ę�x�v��B�ۦ��a{[��t���|�اl+2K>kxJ�ԍZ�ʍ¼T=����
���1Yq4�"�?��i8RgW�C�������;0󽧿?99��ӻs��-[�g/M��� ]�g�v�P������T ����Hi||w&������� Ө�oS�=5weIF�M����gOw�S�D�_&�\�������ՕY�Պ	�iF�F`��>B�����Z�$w����뇇G�Z}>=�C'�������u�{hd��;��zfe%
��U�;�+�O$����	0�O�R��p�Ec1���|�O>��`��h�L���y�ש�����6��������q�G���m[6f�v��iA幎*�^)^r��
7��Q	�o���o��out�����h�����>�C�y��k]�;���_rmV��R��ѣ�����Z�u�LZ [h����m|�2�c�]t�+CT)pF>g�`�W�P�05�˒�_]���&b�3>lJ�s��hb)�r���P*cMM���DZ�\�����_�=����w+UK0��G�_#�$>�)^���� 4�f��<�Du��n'��`�Б�
�)�8.ɯ�g�g�?~�7b6�*���k���p� l��%\�O�Pnsr���X*M#u;�~ǵ�\��3�X�q�x��ٳ¼$G���!R�ã��0fp���yf�m���܋+�s �C���3ƌ����j`�_�4��ӱ du��US�#⵲�DN'�Ug#M�xႯ��ڞ=�>��>JϫטǙ�P����Yˍ�J&�w�y��=��.�������SL��4�aՄ���$�f�P!���� Ne� ���Z�-��_�Y�ju��"E �Y+��x�Iޡ�
&�X,恢!�gβ�
\�LSY7��qڕ�ި��u�O��B@�ܹs� DNUi5��LCh���mː�������2��]���o��V<8޼���3ws�`�	���KdP�� d��ʴZ �� N����R�TG�^�0BRJ�hD�*6}9�
��N�I�AB�t�h� ���C����2uV["�ig�h�gcm�9q�$��[o�Ɠ�zS�>4���R�ذ�d��{�%��'0$l׮]7�p.!�b<,=WA��(� ��T0	�w�`~����8��'�����qb0��e�s ��aF��������G���+㗸���-B1��:�k�V���cM��t���O<,'�mNĽ�>)��/�L�"�xp<�K/��va�
4[��g�dQ%��� �-�]�*�s<�WC����G�0`ؠ(޳M��r�	��6�<`���>0�L����]��@sL�!ǰ��`�����Mu�3�\7�Z5B>���j���I�ԄȕLvK���9&��o6��w"9�b@���bz����>b'e1`lLO¡3"x\���9�͒�r+�(G�4�ofm5�1y��+9!�R3��F�Z��.}Lt��T,V�F���޽{K�JfyW��T�\�#�f{�#���`�Rp����܅��r������[������<
�r��K}�[0U9w�]�|k���0��4�r���B�-�B���?V���5"􏱂~�I�h�c[vSS�T8t��k>q�]]=�O�}��'��ybǮ�7�tSWO7�
�� j��������#)y�d'�2����^6���퉙ًg&��Цͽ����v�k�����g���ض�]�Do(�uw�}�Ώ�2ˏ?AN�/�����i�C�-�_��(�)���I�;o��C{v���r2�������.����t�w����3�UǷi�v��	�,�%��������3b��	�Ǳ+8����(�M7��4���N¶����ۮ�暛o����R�L���뮻����۱c)���M��������jɀX�D� V(��P�WB�( ����}�x�V��g�=y�ط��O�C-�f�;���^����>�L�k �U0���h����e?1"���{h����E�v�39W�j|�,�״cKW.q�C�#Q�ɡ�۪<hKn������.�PY8]D������%ܗ;�ꖎ
��QcJ�ف8�@��%5�h+����̗���*�Z�S���T�T��� 4ǷocJ����F��	KuA��!Ļ��o�Ư (�K3�����0!�QGC�n�S�`T��"�����jP���ڒ�z��]��N��,2�`#��ƌ�����s04�_���l<��;;���I��[�>�lsiT���+�\�k��}]���@-~��_=rt  ��C��u������@x�$�C�X���XOQ0�x�ťՀ"qՔ�x��
����E���8�'��8q���{��׿��#�N)bcZ�b�Л��Z(Ƴo۶m����]L/B �ހE�F��2D������6hV��!�T�}�.�<�/�\��i�&����^9)�[;<?�g�ߍ�`��Tk'rt�>w��L�d��r�e޿"��������ёQ#j,�/pl
wO�;0h\���_����{��I�h�k���+9Vj�֭�H�[�d����I�2c��W�h9��7Ţ8�t��x|BL`�G��2P��m\�n�T@"�|&&&0(dܚZ3���\h��xp̓�� 6�s8��#�lɳO2L+�	�j�޾V��r�뵈Ooi�V,��;v�5²�R��L�P�8��O�\;w��P�y�
��9����Yȁ;� �D%WgSf�lN�g��6> �V�Gãq7!ǴK�X�(P˄���HDW��l4���l��K�@����E�������!8�����t��^��\��ggۘ)a�αٱ^<�Ls�P9|��J��ׂ̄�yhX\L�"c (	�ׁjmr�KX^�O*�JWۢ>�������'�H��+C,� ���<'��t)F���ṘA��7}���$R����4��X2�1ۑ,��>&\�R�Cc�y �v��矧�z��ٳ��U܋z�֛�<G�M3ڒg���0�~�ur���ڇ�lE�q�?���*'#1�7wE�� �jº�}́S|��3F����I�lZץ��y���f�}���Ă~�b�P8`4��n@q!���CW�pa��ǿ��s��p������#Т��,f8k8�������YAk44U3E�o�X�e@ [�֟�PtxhK���V;���������-�O��0<4���7�z2�����ٵSg^ņe !2t��w��d�W�����w����{�8��(�j�oa��|���S���o�+���4��+�B���<>9yy��=��p8v�_^�T��-� P�O�lnWU 4�E�*�d,&`$˾�o��j��+��$�Tq8��э����8��m鎱ͣ�O�1}i�GL�Byk��L�2���w�/���F�u��O���o/~mi1������2�penvn��^pݩ��&g/�A,:;;
���$%�?�̓�-Y�L)�4�d�oK���9��1���*������ u�zP�7�xc��#���р~gǕB�C��T(��
E|�G�I�W%�����������?0���;�[	_�㉔O24`a�ʓO<��˯�mP�(R�|�ޡ���l3�[���۲�.a��&%i����t[J7t���v�ɆE�N���X<M$�!�0�z{���d���U�\�`�EbQ�m��dV^<r�U��i;�x���WZ�f-��	�*uo�f�7�|��^���"E��������ݲ��x�C�D흽�`h`h`hh0�r�"p|O���e(�ҖJ,^��ꗾ|��9�6��`�x��fDW
�Am���o߱{߾&�,�Z��S��~�r��~U+UK�|��.��D�`	����� �1<rggW�0J�/ ~��J*�Ǟz���ַ���ʹW�Eɐ��jeiet��C�k�*n�Xn�
Й�EP���8++����t��m"�@��P4@NP¼��د_���?��<�`�R��`;Sg{�A[�)`��%�2� mc��VV2�*���"Q����F$W3ä�P�p$�7j�eb[w�w��s4_�1*�OD�L�hw�8aݏ{�?���zea+K&��3��|~  �3��-�<�,����6י��m'��յ���
��t�Zr�G^XP�Tt��#�<�����!��4�J!,g4:{��~�ǽT�8U��%Qŧ$���.^ś�;wU+�J��A��{٥l��� \��Ŝ(��)�lKc��
ڵk�*l�Jގ���z��G���+�zL䢓5[tC�d״]��p$\*z��v��K&
��C�_�M��a�r��7TM�7�xT�P��ֲ��D'�%�	[�n�N��5��:�1���ү��G�a���]jB�N�OGB��k�uv�
� ��T��c�Z�]�'W�5W�czcye�J�=Q��,��hP*����7\���ԚLMNq�Z㡇~��W�d�1�J�I]r��ՠ��'U�|��Caa P��*i�Zh�`��f����eL�e��/ O�vs@>��y��C�bf����l݊�Vk�
��їx�A&9��M��2L�d��H�HTٻw�:�Y��f�N�p��X.P�t:�(_�78�S�U(=,����3�m�;p͎�;��92<ʾ�P0�/z�!x�zd<��	���]���-c�Ƕl�)�ڏ}�R͒ ��Ӳu�ԭ�i��jy5�۰*�_;��`_�U�l�%��������ª����Ϟ?[oԹ�����Li�mR}�o��}[7o�grT�X(`qM!��*bI�BѦƻq,46T�H�,�riyy�co�/,`��@�¶�Bm�t2��DA< �4��0\��<��l&6$�L�8��ښ";D/&���$��B���`^3ǣGa�ə͆�(����h«K����L�H�k�n��:LlH0�
��f���g����Q{��f������<���,xD��ʝ�O�+�g���q0%�������*�������p$~Ǉ?|���Zuyi�`�����(>�uԼ2r�W�嫴���\ᮗY��m"k�܀���.��/���������W�ٕ���|$�2>�+���uv�+�ӧO�٦A�PI�L}T7�2� (jp�]w�
|��g�}����-fC��"���r2���O~�����w�2�N��?y��E�)�7�ܹo;�\�(���H+XH$��D+�o~B�<5�-~HNT� FX�\-W�}���]]��_V}/}���R+�B��c�@*���={vG���������g_�I����Ҵ|�W�;Ա�_mꋋ+��Ʒ���)E�&N���ǾC�]*�KJ���{������h9���=�^�������"U��.�2Wf��ʇ!	�c���=@��k�~����Ц��ήh�01Y�t�����4�2Y-�~��O~���+���\�[5�>I���J��mpp`ll�j<`�|�u�TG��)U��l�%�`^���cx�	G�����Pgg�B�T6NCǵpM�e#���g|����9�!��8E�٢E�����H�R �t�߾c�}�|ann�*IqI0;�`���߿k�A}` ���ĒO��9�����
�󓉙0�C�Ο;�6we�hHt�\8�T�M���k[�7�©y�Ё�ёյ50`�6��;;��i��� L�Xldd��*�`&��==���Cq�!�PG��{z{��a�(����CG�??��C���T�ݷvSm9&l��f�]�wvuvU�eLECD-�T���X/"�J�~���<���?�<i��9ĮJv`�j���p �cǎcns�;���3F�y2��;vl߾G8w�h5)�Aj	�ʶ�w�s#���T{"�$(��a:�P}}}=��Mb�U;;�WWW�z���?\(��I.��,F��F8Q�������%��IV�6UZ.���V�Uɂ�5�l�+U�v���K��7��b��gA|�AP�������=���L���c�Xw���Be�p��O]��#�0�;�sssLS�A����T�
m�e���4��.��������:��<����}V �w@ȭ;a�n����TJ�N"O)U�RU�w�� ˸r<��2�����������1E�8;��'S���~�� ����,Lx+_��q�__ww��mۉ"���`�� ���H��e�/�R8�B��@��Vŧ0<�pOO���0�Dc�X��G����1��/2]�G�Mq]��R�t/b.QU�*��w�|�c�2P��icE�q���`����O*G!8���F0W�$�d�r�����׾>1qn=��f(K(_��G�����/��g�zO%�*}r@SC�j�O��񏦩N	~�z�Vmʾ@(K&�\/ĭ�pSL��2Q;��uב�S�ɧ�|��83VD�Z�蠵�M�x7�p����n�Q'��R�ش�h�� �o���+�ġ惐���E�Ѥ��ӹCnm�ŋy/������o}���89�m3ۤˢ�J�xt`�������Cf���B���&_�U���"�Gd}�~��U�65�Pb�x$�=���2A��(Ŕ�9��q�ĉ|����B~4	c�-����ρ&��
��� ���P�4�z�{f0���Č1)"S;�f����)jJ�b7�r�p(\M�<+�?
�NRM~����_#>5G־=;~�S��������M���[�T`<�� >A�7�:��WOxW{�,�*k�ܢC/H��^\Zj� Fb�˫0۰�1I��7܏����U\Ǻ27{��eR�n+s�����M��d�����={�7C�g�9z��z;0��^*
�ԧq��m�D��+�j/]���
e��u��;p��#>3=M����=�6-8��'g��zaS�\��'>r�P�`qyi�ܹޞ���M�Ht���]^Y2-R7X䠪��FM�t��7�x�c�@�z���7�8u'�n�O״����/6��e+����������ےmF�x���~��VXCUm��^Dᾗ!�|�?%��$H��@����fs�L�r��c�!�R5���+������Z�\(�c#����l���D�xH g:<3��zݨW��6������χ�D�F}�e��J,mTh%�׵E����r3���WJT�Y.�HgW���E��>(�ޑL��������J%�lۼy��Yˢ#3
�zC�8bC����o���w�،�w���۪Պ ,rU�j[D�@O�%���aD��NK�2N\�=�Jaؘ��{� �̍�mN�ۡ��ܲekwO���x�����'��f������#���Ï<��7���O�E�Q��A����O���SS�t�?�A�So>��U;DƍC�{a�n`�T[�=��?����;���	���S4^�!��b)�L���ث����#�fVs�HD�:��b��1_ȧ��`|�U�\*���Ȉ�DD����	fw�vP8�; n�� ��~���% ]���w��җ�nm-/�.9�[��i��i��={��^���� FPUlm5���l����a�cikKwvv��: �a��`���~�#�H@D�Ǭ`>��cG�����ӟ_���ʘ���y�b��w��
�NITf:x0��^�F>Ae�<D�\*Is���������zu ����v�nIJ�k ����m:>��p���˿|��12ul7���*�؁�*������ �@v� ��4�K ���!�x���8��%��6A��J ŭ[�q;;����cԬ�����}�Y��gE� t*�P�[�I�s������C�]˶}[{�P,@z�5h$5L)�a�z�F!�x4`�ΎNѲ�P`ut�C<b�(�M�d�V���|��_~���E�7�nU�+"Մ�(ˢ���
�684�h���Z\\����l��6E��X,�#� �� �m,����?0��ёJ��g�X)��o	t����y�^���)�����7j�Z�7^ɵ�	t]Y[�n�ިך�H'u��kԍ��R��S�M�� �޴i�8���0��J����z�o��o��<�h�dAvE3#.;��z�Vaq]{����~ݰ��$@���5�f�R/拎-��) �)�H8����������n(���a >�(<�r�յ�������_�җ����F[�m���B����V*Wa�C����Ae��R  �*p$�(-,-es�z��jK��@Ec�b[�I�**v$
�A3a���w�ܼe�?�o��o<���#��vm��;�`S�u�ɵ!�[��5����yQ(�3��~t-���Y����hSw`[C^� ��V��W$���n�fOB�����Hp�j� v�r&���8M޵��x���+c"��qz�(�kQ�ܕ�P�70K"��`��W��}l1�;G�����԰��(�(_N0�kY�4~&���J��[q�e�!W:q�'?q�'>�/V�.]y��k�����ue~QQ[�l�&��q���"l�Zn3`߅�0��VrK�ӡh�Ҵd8_(���kvmVCa&np��q��7j��_����P-$�$95`�޽�}�z+v�Ay	�bʲ�Pww7�A�"�fn�̉�0��^s�����]��r� 7("��Y;��{��X�F��5Kf�Ay��������]w]<��~ǭ7�<s�n4��"Y�*�*��)72�>{�f��O�*~�9��Y��Nl�2�R_�@4cgR@���#�9��N��f�������6�j�_n�K��7���?��?��?��`�|�	���~\\\�� ��h$i�N�P�J$��Q\��i���S��%)�@uu��Gy�'��d�{��v�9��D���z�\���7~�7p��=uRD�5ꭞ�c̢'�P5�*�I���~Xt�FF������� 8HKN&�i7kM=IU�ſ���>��0�A�im�)|R��z���}��T�0�@��h|���w���G?��~� w���$��ٙ�vr�B��� �	:���ck��!�WR�-"�L���o��O<E����f������<'��P۔�|>�����K�y�_��_r %�(*]p�`>4�1�a<���V�/b���I��\�DJdz�P��^�͆�X++�Ǐ�ZY�M�=]/"�$���$�������ȝ��5A�P�5�g w`]�>}�{h�+�1�!��$z������Y����٣'�|��_�ƕ+�BQ`O�u޵Ҵ\���}镯~������V�Z����ҭJ��% Fܶ}�9��cMM�-�cH���
,	����M�P)���`��_?q�$ t8D���t"���[dE��kO?���w�=4<��
|�	����$[��4�)c�mI&tJ����"^�P�>�rI=��0����;:0�o~󛯽�'5AtqA�~��TN�� ��=��=�ܳu�6�p\��t���4`�P�I<%KK+D:���M>,�bc#%yLq���G���=�1|A?H$r�����կ�m�z�-��LM�?�l�a��tFU���;-Zm"aSE[X(p<n��l`��+����Wa�a?r��G� �~��ֵm�򥹩�)nд���hs�XgW��-+�[f��u+L�4�*ۖkZ��D5�Uv�EKS%����&닇C�1Q��cE��� �AnWhN��#/}�����g?I�De�Aݥ��؁ue �:2:T���<��z��Cǜ�{���d��t�?5�>u�����	��`���VdձE�8�rm�E��J�~���W_}����⧛J$��T��-+�D�ōz��bb~򥕨(�a���K����7����"/T�W��?Qg�j���;;�-S/dsX3��c�=���@�yF͠}*T({��g< n!�[:pv����UZTE�J���n�q[Ƿq�R4{镗_8�"��0Vf�o�x�r�	�Z�U^}����۔h�-�B.�Y^)Uʆ^��	�5Ksq���ħ�1������i�'�ݝX�1=�.l�R�<q�B��x�JQ� �b��T��ӣ�X��9��`�~�Mg"{�6��H$fYN6��$1A�#s���ޛG�Q^������^Y���҂$@��,6k��ݦ���y3}Λ7��9o�������w��v����6��`��1�������R�����{fdF��~7�S�!�%$�Ns�U���/�����~��������?�/g�TT�OR��E��eQ�RPt��<�.��ic�[//�*o����}N�����O�&FFF0���o�&���J�q'�4�p}�J��}�W�����������޳���}�
��]	��b��?������^x�WE�s�r�?���E�v����o�s��H�>ݬ�#������p#4���q��FG��?�	&o��?��kO/L�L�@�C5rt��6�'.Z�S�|�&�KXc���������Gr�|G[GOo%y��_��L*g�%.m�e|�3�oټ�w:v��?|tb| ޴k�N	b/jP
�iV7m��_�����-.�V����೿��i�Й�;N�W�"kx��84��v�!��U�&(
�����[������qŋ�F4Je�͈$��FG`��D�%����wS�����g {CU����~��\:�5�l��ޱp�A�q��Fw!�����m��R3�P۪���@�E�����'��:��׭�ݶmۺޞ˷l���z�H�ZkX���B�.�\.��?}��G܆Z���Rev*�@�j�e����F]��)�0>6
�?u�u	h\�&���Y��;B[ �a0�_~9�O������0-� ��Ru7%���۳�+_���={�r���ڵ� /S�y��CP�h�`�i�PB����䧮�TϚ褀��*�{J�Xb$XA�(7������A���������"�&�����e 	H�~��g?{���UM8��O�sQ%��#���R��-[���Ǵ{LG$r[��;pn)�E8,��8����-� .�a�c��zz`�}��{��կ(�Ey�$�[�����3��s�}w�y'f`rr��T5(�W�z�Aq�H��)����Q<,(�О������lA*���	i��o��Z�5��o���q19c,����ۮ��5kצ��DN�����m4���0���}~��ɉ�x�	�0�d2���]��7��Z�ʺ�{�§R1��\,���q~Z���n¨����;�� !�&r2��Qc$�]�ӳ��#꼚Y'�����NE I��58���g����O��رc�e��W���t|���,��)�����?���2���,�)�	c$������I���w���ת&7B�nf"���ĳ�'��/_�=/�$S��D���@}̪���\��+�����>�Ғ����T�)-�c0�;P�J�\�����!�`~��)ZZ���#���#������~Αk�cb'˕��j\��Y-�C�7nܰ�2��<E�-��G&�+K����H��0*ޠSn��\̟)�-8��\Nw+��׿���^$���F6��.J~]
ёP��W������ݮJ���f�jc-����2��{M�������7o�
��BSni��m߾{��6oذ��{�IO>�&��Xz��*���`&�a�����n�[0Q0G�'�T�^��A1l�I)oD�7�I0�y��g������꫹6�����o����<3�Ú�'\kMMUISCC�P�lӥ��X�T,ٔ@Q���2��T�p�Y�������)D�P���LJ�}����{��޽�!�R��|��1��Y��E��j(|��|IP%tBq�c��ۚ��e��8�ħܣ���Ɔ��R���J��K-/�,v~�u���>{�m��\�?0�����;x�ګ���?�'gdhd�-[.����U��[�	��F#M^@����֩�9�^=��t�|>%��s3����_*d]�L���������+���B��^{�&�2,�N� ~��/|��M��om���T+cC#�>8:�������L��t�h�$�x��B�Ti����Bօ7�_�3(���j3R��8�����7l��w@�]G�BRoj2rth�-[.���O>�0����>Q���ȱ(���9��:����������W���m�T�������jͪ�O����^ʙS�X�\tC�Ixe´"�j:�q^���6m��.�	�B���j����M�vui�D"�֖$�a��	���
aZ��� Z+U�'���=ã�؁&�ݨ�*=����80@X����	SS3��߾m��٠��P�FU�M�z�-CKb�捗m���ъ�R�ֽ^56���7���O~��{����쟎��\=ss��gPʖ��Dj�P�z)𛙝�l q�B�3�5A��H��s�
�	�j����`�Y�`f`��c\n��7���W���W_��Lr{6nZ?>1�Q���CC��������B�^s�5ݝ]�&���4[U�vO"OՀY��c�xWWw,�uH7��"����UR�b����G��9��\5���V���Q�<�C�HƳ�&������R@��3S����|�LiR��&1H\��k��b�����'�x���~��r1�RǒS�q�7����~�z����t*5<8T܃��� p��K����8`�vzk+�x�> ��xk�4��?�ķ����T�O�if�-�ږ8��7��(�0B��G2�O]wlK�S��@�@�L��E���N ��w$"��ԉ���0Q�v�뮻����	s�Τ���+ ~3��>��v��<%����9L_�=L8;��;Q�$����&2�\���e��[-��5'��@(p�����W�������_��M����A�ՖX���	DE+�F���}��8�����X������	ǼQ���i����`�������\�90��8� !�kn�X_�?W]ye��� Cs�E��� 4�,��#�'(��r)�l���7��ఔ+�kcƨ  1���/?��slz�ߔy5��K#ۃr�xo� ޟ�����[.�ꅭ[� �V��z��/�U��d�!�Z-�a�@�����8ꂃ/j<\0��������������H��:�P%��5B��K��F�0������CC�xx�Ƶ�` ӕMg[�QZ�Ly\tTA:3;5;��Q r�]��X�[�=����ـ��y��'a��3�"W7	��*+)N��"6M�K$y���M_s�5����)*>a��,

��0��>N�� B�x���)���%Xe�<��'��t��d�.�z���4�ON��v$[��c�X���,�
��D���A�h����"hnn����b�v��8k\��Q���ￏ��C�{��e��-W*���.]����g��vk+�<::�qa7�`�9Y�?'''���D]� E�t�˟� d���@�:�����_����Yr!L8N��vŖ;��s������b����/�����ز�rW�&��~���E��`j��`������8~� ;b�(_ȿ����������]0�����ãͤ�S� iA�ںu�E3�^�����w�Z1[ڪf\���[n��gmW �cB�����y���d4���JUw])�U�69K�ɾ��P��T��fQ`�mYX.D[N���`WG���n��s���l����"�W�W=^pIw�h r	E"�ãc�*YƔI��xa�j�Eu�7���m_��N�O�T��j�����ۗv�M�&Us�r��A�����H��b�L�`�(Z�} �X�~���??��t����wmh���Ě���d��'���IdP�[����D�}�\3͟=����H�I��j*�ՅG�xj�t�B��| ������0���v�ܹ��k���M��X7�� ���C���q���^j&Q��f��p4�KQ&&G��W=�c���*�Ü��[�199͉T�D��:Uڸ��5%:���Bj~~dd
t���`�MN�C����]׻a}_ooϺuk7o�,�A�q������TXA�b��MɁ�|!��z�w�y��g�ű�`�������c��U�D��/��c{�Yp�
��������J�E��r��yR��mcф���c��P�n� 
���t����+:P������O�|���"���M�`3^o/�W��f���?�^X�,ttvp�gaɚ{�E�#!,��E�L#<���i|<���Ǟy��hvȍ�RJcn|5WJ��Ͽ������ՙ�L:C5߰yGH ��� xkk3�+��~��>�=?���1�O=��7����I�9�/��F��� b�=����Tժ�ծ+�Ϸ��}���m��
�e�\�#zC��
���b%��R$S�DB\T���qeX�`r|�k_{镗E��2m0T��\>���K��(MҤ\.�Er���Ç�r�n�Dȭ��y�C�\�OQ�_w��i���V��ݰZ1� y:\T�GE_����o�[?�я�&�p7�a�� "���l1�0�.�f�c�������_�_J\5X�u���A�F��9&�/��Fa9��Ȉ�8�8;�߿cǎǟ�Q]�nH�q-	�S�;����L���'�C.m��A�X6���K-��O(�c��յ��w-6p2����Bqavv��������`<2�w/�6��`D�A������ѱ��1,���>,�]���5���7>���\G�{�&��`2�2�Cy������>���s�<M"����������zWѥ�;>>948�yZ[�D�R�c,�f�!p�:����W����>��oS__�	�2��A�Q{[[{�A���g�}��_�
�5�N�f�2��Î���׬Bo���%�Үn 
��G3`�2Cf��	��c`3���&=��+�tGG'�鴶q�K��~���@�Ԣ�T�Py��-m�u��{�.�+���Mԣ�x<J���sW�ZWgwK��A_D"��V,V �j>=!DM�� ��I]�������K/��Nvu��T/�;�a����$E�R�iV(SݪC
e2i����>G�P�����pӎS�o�G�P,q�`�D�B�j��O/;w��]����Yg��	��~�x<��}��+����N�SWm���M�����6n��� ��8_u�!i;|�$9p9�)
7ũ�����:����)lZ�2������Qݲ�6n�%Z���b-d
C�#�k���/0ɳ-:���.�Ȇ��Ճ
!�J$~�M�Y��uz��[�g�ӿ~�ŧ��MY�6_�%�Tr�XK'@ �G�VP�6�h3���>���:������Y�B�BI���B���\��2ݯg���}�ٹ_0\�V�6;;_)>^�a�(������ޱ�k����o���n���7}��o���[����}�������;no�h��.����?<Q��h��64�b�gN�sB�
�������f�����.d���
?m�m�]]x�b��%�
��799�*,��� 
�A/��T)L���������ߎ�n��X1a]�g�\��;��Ri�%te�����m���[o��w֯����Fn7�[��J��?�a�R��ҕj��V�Ēo��?
�{��ď��;~x��!]�`�Ay���Ã��R�	�6�R��F�a���z�:�-� FF�8�s���A"�!�)
�=�Wtnb���P,Iv�F�z(Pkvvf���_��3�뚡�?�W0����CT��"uGĩ�Y��0�§h�ݻw```ÆX#|���l%[:B��G��,��x�­N&-,�|������'��@�ڽX~�[PU����ɜ��ˢ�v,��NLNr}1��������ؐ>�$\�Dy�Ǽ>�C~�������)�~��r���f?�J�ͦ>�ފ`C����{a!�k׻�B�-�5t�u��B��a׵�������Nꩽc<L%�}���O~r�}=6Xe��'O��+%�`3� V�	�;0P!�H7\�l�j�a��������۶m���	�B�s"���#��I�vF�{b*6_���a"����{a����T3k�'��T��__q:�9� �v*���=vSs��|������qk�d������k{�9��`�F�A�~Jc�,8���w��G��^M���NuZT�OJvJ%�U`�S���={�=ڷn�ؓ��������D��HT�0��@0���gs~���|�+�=�x4�	�P�\��f��*���7	b׽=�����~��߸qcOєg�i��qY���� +>�A��]�����k80����h4���~��MǏ��]w�xx�6� ��9XǓ�#&�!\{5]�x9��քC�ߏ�3 㡽��Kq$rz�ʁB��"�t�H,�/&��ئn~-	��+_�����C��y��Uqz [<L|���~]4,��M|�6�Z��G�=bP?��d,><0�--���1ԦYBVw�w����V�h��dzب��
��_��k_�W o�Af�x�1 ߲���
R�\*�B�ai`lK��GU�U����n\�"۪i�$�AM��������L���U���L�X�>
���=��7������h��VN�gc��vA�,2W�FY�f��66<:?7�v�z{��8[���]��ghn|)��:Hq�Zv!�T�Ss��Ύ|�@�d�:�~�Ν���ҋ�t�ԭ��$fYga��)��2,�����*�+$��G`\��Y�~��� ���<�x͚��Ç��isI!v�֭[�p��#G��Ǜ��N���y)�Y	] Ch}�V��U�����[oř>v���Ç��37��H�������"b#Q3*f��d�x��0䩩����l����?Q��ݝ/��&�Z;r�5=��7B(���LMO��`o�FH]&5�#B�z�7`5Ԓ३�V{K�u7ܸ�S�;�^����C�~��Ó�7oݴ~��m�ƆM۸��%�)������0~���f+cgN!ǄK-��Z�@N�'ʥ��5}����֖�o�y��@�R%`l��]���~���W]k��,;ޞ��-7|ꆛ���;n��37�t���rǟ�v�m��r�����M[�� d���I����O<��'�r�� ��M!��J�qJ�Ҕ=�[{�3�k�Kf�"���YH��`��cG����u��m��m�,C��'�(�0e\&���nm��s����6\�lf�{����{�z�gã~�ʯ
�
U���Q��r1.�}a8"ř[�q@�M�FÂ��ݷz.�^��Χ�����mm-mɄ��j@n]���7೪y�4LíGb1ˬ���K}���}btl����}zz{#�������,��D��g�Զ�n�9jt�9�����={`����L&��\I�#�p��[ZXH�B�T ��`������[��a�?��S_��o:t&�*3�L��A$s�3u�ٍJ�<�Td�Od�����J�*������?��͢�\�^��X*�U��uݎ�}T7��C�ݾ@@s�8ǆ��q˷�~����w�}�e���R�b	*�����Bx��⤣�$�$����=q�?W�C	�Ab�N�۰~�M�:�\-���p$�Jli�$�0���s�����������Ջ%Q�brʠ£P�$>�l�0S����b�7���;q�X,]�v-�0�]*���:��7�ߠ��dK_^����I�Pd��!�1o������z`d\x���8�fV���<���RV��@��T|�>��p�>����~��ֶvm�m'lY�
�ٚL���e�J�h�Tf(��}����ջ�'�~_�?�<���_y�#r��< �T�%�Z[�5��[�!I�r�*�f'�~0q�7�2Q��"�֋��u�'�-01j�JŶ�/�������?}�������P�Z٤,�[�A�>��h�d�s�.搌H�#�����OO���-��� ^��d"Faz����*��)�W��J���S���O<�ow�o��&d;�� �59\�v:�"R<1U(p��0��|���#���^�խL*�f���/Ǌ��utm�[�5����+W���o�����˯����|��_=_��2T�&)��~�C]�ʖ��9rF���sc����y��b���J�f ����뢙����4.*�R�Q���ѨY���y��>�s�F�קh6%E����L�º���F1@�P_ǌY�s����ᡱb����J
FK���hk0���Z�<�?��P�&[y��w���ݏ?����<=��Yc���Ix*�W�3l�o�D]��̚u�x��|j�ڞή��r��|����`V�p~�ǥ�n/N�zA���vy}~l�R�tϽ���/����$�y������!#��ѱ�s��J�|D�~���M2s�����+�&C��e���l!�z4N�Z���X��&�b�X.��3w��������K/����^�i$Lwh0�p>�,Q�6�-i��a�k���q�	���m�~�?��}�R!�I���%b8(c�c{��)�<�J��>�)\����ށMLNr�W�+���<F*$C�3pq���~[�V��	�(�L%�r_�usך��]���S�+����k�C�þ��۸n�U�!�V5&Ք�_��*|�.^Y�bp��m�����|8�CGX�Lf.��޼~����̦��������pj�ZiՈ�Mm�x#6������_dC��W_堼�j�iww����6mޔ����MO�N8t�P���]���ڒ����%:�K�հ8EҎ�;ϬUF��ISE���m�m1@����v�����q3�(s�0222??�����M��I�"���-�CI��˂��%dp����w����?Q��˂M�a
�g��1�de����2O��g���8��A���-9r�����!V��a�D���@��T�LJ�i]�<��3�<������==3m��@%4�T^*��y �5Uɩ�J.�Xh�w�رc�T���߸q��c|H|(�`XAP�����lv׮]O<��'~���v��\E"Wc���433�JS�T)Ӛ_��r/�����Q���ɓ��� p�����}���$�"<4���}�<�ba����G;v<����v>��[A
��FK2�F�����4�/'
m�\ju�p*�N$���/lݺ���ۢ59'�`��e2܆�cĦ���u%
`�����'������SϨ�V���%�cil��g�u��K,��j%5��_�d�=�I���N���H(�L�P��m�+����ME�Z����;w>p�������'�}^wմ�)�{�҅�Τ�@]Xq,�/�_�nݦ�6�	���ƌza���B> +ell��_|dǣ?z�G�E��K�`c�=T��b�p���>cN�a�M�qܹ1{ī;53�k��ٙ|>����N�Eu*��'b�0@����2��	�#�ry�{�}������}�>d�GZ8�����x���Q�j�U�(\?::�{�nj�*��BT��2!�JH%5%1��3\(W*�JU�Qzᇏ>��+�����G\�<�0ϼ:�ޅ��4�d�8Vݜ������cD�9>>�X(�V6�A]�T��B�X��Y����/d_m�#�x����9bV�n�B�5��S済ή�"`��T�����	���m����BQ����������g��h������Y� �g��{�����|��w�G_M��Y��^�gnn~Ϟ=Ǐ���"�4������O���p,,�`z�Rb�a��\6��o}��'�ص{�|��ʭZ�=_+U%�UJ,�Q��.����Ç?�����֟�� �)Y@Ǿ�C��Xn�955�G�`��{�r��Ƙ|����"�\�l~@0��
�4ީ��_�P�\,;r� $p�޻�'�`g؂RE���,���x�P(`�Ŀ@E2�[o��������t�E�gy�%����f�燆���2���Z,�Pq�9LS$����y���r"k�: ��߿Vf)�˱<�d\����2�D}}�֭����w�v;�ϗ
E�\�l*������~�5<��8���oݺ֖�����߽v��Q�:�Iۣ4i{ϣE��"'�'���G)����.5��nO�::[u�17����ԧ�ް��D-��k��q��~��q$T��bZn��{!�]����
Q��ɺE�&%���W���tj����h�h��q+b�u�/}�K�]v��0l��/{2�kj�K��X����'/3�����D6�kikY���5"��%��4Ǿ���}A���ѱi���	Ȕ����M�-�FmXLݦ�s�M� ���ԃ޿���ۿ�߮�b+1ϖ2@��r5� *劅r��_<>=�-@Ǥ&���#?����L�"���L�8X�%|xU%�b�w7�J��5�8$������_~����NӬ�r�-�W�'�%7��ν��z��w���5��wށ�jn>�	�@�b`���^O�v�b����A���W&��ۿ�[.<P���9q�D��k�F`1N�O;v����PN�{���o���b������I��������_%�8PsK`�>|��w�wQ�_#.fJ�9,^�D�4����LLL��S����[UoCL��L��'��fqE�#��aa�QBF�
D�)*ێ;�j������ڠz�XP�7v�8 Qe[ca�Z,W�P�##��'�|��=�흙����\mn��0"�q��� �H�#
���ѣG��4�����XK�ۄ,��-���W���lڴi۶m�	��1?���q�e�E��=+)N��C�o�'N������ٝ_�˿�K�cۆ�+v>`����#���R�PF���}��>��ILI(>��I�jy�����Vkܴ���;r����������[��k�chp �[�&�����r>?1>�&�Ɂa�d/����#G�DEQ)W�� :����XJ���zԊ��B���e~��wCE�Y���7���ݍ�co��VK��e�������?��?v���ǎ��.X���ε&�Lä����T0�0)mQb��<z�x�+/��e˖뮻n���
G16�Mޙh<�]X�i:>F�'O�<q��;�-����B�:gA���j���Ɵ�t�׿~q׮���n�����,b�}]f�|j�B:;4|rp�dŬ�g҇�{���@��"����PТĎU�U(���{o�k/�p��Wo߾�<F���kUS��߈/Ѯ[����$m^���;w;9 #�����E�SW�]Nyx����tbY0)���?�?�������+�����E]�=��|���M�-�e���\��P(�$,/r�P�:gU�,�A!�YX���9 NX�o��6��x��7wv���5G��9�7��2�N����G |~���dU/<3�0� 7w^,��k��@AT����S��b���tcC�Vżhxꃴ�F;�ڒ�ش��P��@L�`.W�Q)RVa��2@�$�H�6�����VE�.����)���JL~����7�0�VHiAKw>I���W�T�~�E�t�j�w��n�;]#��5�HP̡���J�����j5+�'�-�\Z��[≭�_��̦��R�t��'���xCAR�8�)�����c�+�9 M�u���)�,_+�
�J� �A�[��hk2&�V.YCH�B�� !&ܪ����ՙ4QC.����p��qS����T�W�c2��SO�����^{5�b(�.drUAQ�W,U������t��/yu����/��W�.��eu1A��ҥk9����u���� �S�!��� ߣ��|j����Ǣa��p$D�P:�}�}��sE(�T*���0�atWTL����G��2�y�r��>N}�D!�O�S�e
�=�p(��������nn6�(��轣�QU���cO
����4x��M uѷ7��#�F#��-�9t�s�=���^��ørfz��O��駟�ڡ����٩��\�P�T
�J $�\�	�\I��ff�D��"y�����,�-��Sʪ�[�=��������_�_���O�s�=@�_����^��D3�2�d�����O�
�>� .5}䧢?�i�پ�-� �x7wk�b��?7?���u��˯�x�+�؂Uÿb92�À��~��S�|�B)_�* ��Ç�
5���M���U�U_x�{�w!K�X z�Q��hW9�.M�z|0T�D���_ؖD�mF�4��%�l��C�T��(W���C'w���;��n�����-��ԴJ�����+���/p[�摣':��/ ��|�9�3q �l��A��}�Y���B Q�0~}.�I���ֻ����;�w�H2&������E��j�/����?nV�VM�L��W�Z����ب��������a0�V���,x��]���={�����N�3��뮻�eP�L}rl��{�;x��6�{��ǚ
cU�Uݰ�=��L����ս��R��������"��i7\�?��?$Z�K��/��Ǵ����\�853Cu&1v@��؋ɵ�'<��G�������4��8���ҿ|�/��24���/�<��&5���:������-T(�lU�0VK��R�q�VXE�9l�J]�{w,�ȗ�ө���o��;�����hKn޲�r�47㣏>��C1�7��w)��+���G�"E�RmT�	�L����D=B)�L�C�K�6���B�s'�B�ӟ��7^���۞h�E?.ڮ��@�n�����w�م-�o�>����KM�񮔣��J��U��R���C�'O��]�鲭�U��~F�-���ޡ:!pơј�R�_	ޜ�u��"'������>� �*M�
�'�P,A�b�A��K�}[;�u|�yN�%���+]M���O�v�S��<�^�N�=�Q���*F�gR�0�-���.V7γ�@J�l�A��Љə��֞�:�p*�`֭
y����R�:P�h ;ªI�:=�[���W�qV��^�hy܆&Z��������d'%��W$�E��fӚ���)��v]��5�0��[���U�����5:!��T��Nt��.x�8�$�-d>���'�^��i!�n�RM7T���5�m��Ш��/�݆�f����ڥi-k��]�|�3��-��`�>�`qfj��+/�% �֛�&&;fs��\�[�#��U!�Gs�u��%p��H�H���3��LP��|��'w���mW���������W_}u�ۻ�U ��Fm����~��Ev3�Me�9����+���$F]�$��koK�^1'����1�6l߾����sύ�N��Ɖ��D���hG=�(��� ���L&]��������fd�"�aQ������g����3������װ��g�=���?I#����
;O���Y���7y̎�4֑;d�)�I=��jހ�z�p��G{��X7n�Ȝ�3P>�:r�X]x�)��b&&�*�D��jk���y3o�zrh����gn�	ߒH$������;o�=>:Z1q�9|�t���\��A�D��.f��	I����l6��yq��[mZ��3SUOܬV�Ɂ�t��T:�Ҕ�n��VDÙ��_���;y;�zP��W�]5MYmO
q�F����4Uut��E͎D�E@*�3�������8+B (o���e�c�sss�����������l���8^����~( ؓ�=���ꦄ�����nOŬ:t��ѣ�d~���7o�(�S_c�;Ｕ�-޶2��&JɫfM1k*��$�j�s��f�4��Ѣ�wL99)�נ�\�8?;_,Ug��>����s�3kE�P}啗�y��[�}��p8�m��7%��*�w��T����l��jD��� U@��raxd����+��t��,r�Je�2���B�Z(0�|�	Ί�G�}.tr�v8O��mx}"�-��[vfr|r�{���v%E�F��_br��1��
Q�/\����]"�R�:UiI�����H��d�%
:�^r�y��l�����=��S?�	���#�f�8}B�T`l�J:r�8���d/�R�Ba��]��`������08!`���AF㡣�?<z\W��m>�������i!����o��7������5p�f�8��ͮB�sۥR��6�.
����_ggg�󹗍�Q.�cM[q6G��{~q��?I���E�δH$D�!�h:C�mmԊb?#j{����Sqʥ��,�z��!$��L�233Ch!���/�Y(�͙�9�Jꞹm����f�2R.ܦ�B��PK`t��  ��K���*�C�X�C�D��[!o֪��~i�B��W�}�2S�R��U��uC~����.����'^�r"]sY*�A�Z͊���M��L��m��И�A�R훭A�(J7y��R�)L� 5S�׉Y��K��:�,2^ɨ�}��l���fy�-��3��믿�曯G���=???59G��(@�Y��n$�zH���5EKB]�7h�s�X\���ۻv�Zf������ao`�>/�f@��n�v�ŏ�D��D�Vq.5-\����R��z�I�h5�B�"=��G�JϲiӦk��flll���y����~������m2"SBv�&���.Xc��-X��q�u`;��(����tWM�5�I���g�)��Y9�ۆ���;��BKh8w�N��G��p��>�5Q	G«�}��P�2"'6Ώ/Hǅ����~�?ǪE�B!�^��>Z0L��U�T�h���\��+#u �*����ꥅ��c`����<�0vE8LDd�_8t�&U��ڦp���Z���f���E#Z�E�r��`�3� ��b��#~�}ȝ�3�,��W!6y����?�1&c͚5����û��C,��SG#Z�\`Q	���%��5˲�m�ٱt�i �'Pf��Z���%>�-���+rq[�@���C8p@U]����'NNL�`��M\�NU�U9�������܈@��\����6�b�h�OT��(۾~����k��U�s��'X;�:�fy�b�f�{�+瞂���R�˺���˵2��R�g@zT��3��7��"�C��������U}~�f��>��/Gdϫ��4R�<�":"uK�U"�K�P,���jR��[Y�e1D  ��x)��\Ƴ���di�du���s��&��4�n��I�u[��@��U�a����'?}񕗱Q5#�o߾���f��ݹ\[��N���=�X��"2��z`p�U�*E<�d�D��<n�����:��HͲ����qc%fQ7-���D���0)�[�E�j���K��Ejt��dH^LN�X4)�����@���^*���سg60��{��B�<S.1��c�A�T�ґ�����.�+�v�e%y��+��*cuܢÇ�Y�pr2��1<p& �z�T>�v�j[�9��@(l�����{���P5�^��B��/�F�PO�eV�H4K��T.�J���[sC�M�ܪ[��5�<�c%���.XR'Q�EN�Cs���	��A�N��9@�����%�]^%;�j^�Ks�I+��p*Y9؋�H�(��%�j]J���],l�,�k�R�z��*l �����T�Ԟ�"@(� �]):dZ�_�]�|b����a�I[�vȟK���c�8�)��'Ǳ 5�~�t:�����Df(	d��B��Kg���(�f�s*
��k"D����b}��ѱa���#G�LLL��V�j�R�T������"P�#�x��@>c�j3�<��g�Q�fd��:%��%��'*mhh3	Gȑl����|1W�8���:�z<��mV/��ց`ڨ��ͥV��̲�x�����E���م_���au����N+S����P����a�j6���k� �#F�.�ˤ��'�L)��
�{c�[��0x����m~S��S�Oǻ���abd��ߔVP�5��JJ�69�Kj�ż��+d���+5��&�Po̰��B9nu�4.�
�m�M+��4*7�ǭ�Op֙�̤�������8�>8�YP���T����>P�ej!������W�����)IF�YԮD���;ҁ�K�����J3S��Ɇ��L�9�8��xv)cPN���961=���e�](D���\�Y���ǔ���&���s��&��q��,$�EM����XS����Ʀf�z�ٚ8.7Z[��+U��`�`���"#��+��D�i���u�C܆�S*�!G����~�[�^�I`_�?�CW(��ы�;_q`�͒U�C�r���Ե�T�!|����k���
vG^"o��x��`�.�U����aՙI� ���K+[A���~��;�*�F�a�[�4��T�����Ʀf��ƗT�m��n
|O{X4��� ����`���:h�:vN.��a0c7�d`0�� �1����a.�q�S�7��a�Vɕ``d��aahDa�:B��8!�R)�J)M�n+' � w��R-+"��6�d��k[t��Jｷ�����iHLk�\!+b�7MRE�N4��:�3�a5�	*�hyD6x�A)I=�1��B�rTg+���J��!}�Л��l�|!r�>�5B���a�4���A�j.�J�׵�����A᧨�\���.�T�Ko�n�,��)Т�����\jR��6�+��R:�u�$a�Qn96�`"q����P�� �B΢%[6 ��~/�\��okO֩�Y	-Ov�ǡ�U�'i�jH�Ȩ!�J)�z6�Kݐ].�11B�[��Sa�HF>cժ��b�S�Or�1�+�Y�#�X�Z�}֬��E�7@%�j�j�E�rb�'�)��L��qp��pfM�L,��J�(�L	�5��L�T)b_Q��Z: �
��p
�#F�ok׮ŗ?~6FKR�f�a~��5�&2XE3�Cu�4�|>����V�e'��y8iAEC*i�j��C+����:;;1l���z�0��[��+nݜ�� MnI&���?��Z3o���D.�`���ؐ\��s�T� ������6<���$��h+��$������J03�S9U��]	J�F�@Uu	�qm�ݫ�n'�����g\�`-sֻ#�x��6��TY�s9�R碓���7�����):C�K�8���Y�9A��Q�ߟ�簩�0�x5�"��el����Ǡ4,.?�,�`w;TqC���68p�������D�Z(��	9^������!�jfv��	��E��U��F{�of������Z1~��S��яKm��ר�B�\�'�o+�8|�Dv>���U��I0�S{+�Êቂ��9� �s��
O*?�M�咰s|���nؚ�j]'�H����(�B��9�P>���`eX��w$�fA;��w�IYԊ���,PȹH0�1�\*0�4��N��(� S!�#)2���*=��ƴ���v�����ac�J���mZ"zdq�vrMTc����U���rACb�`wH v�*A�G�����n�� �+TjK>�,X�l�ר���HF�S�����)�O�u�������� �^��f6�
�����U�rpw� 4rEg�
�Vp�G����L$Ya\C{��#�fW�&{��@�$�����ldx�k�!�� �4rӤ��V��4%�.s��r�H�TN/�8#�%��
Fh��Uy{K�+���58�#�r��~v5C��hYD�����$��up��C���X|�R
}�P �hP4�h-A�D9�ҿ�((n�s�b֔hK�:g)���x.��i���R�P6E1��F�hU���/�"s}\��3E��(�P�V,rmZD�
L~�\�N�Ӹ���%�`�����^���	��F�x �U�C��*��]-��[Z��h�hߴ��5݉d����'4�K���M�X*��Jζ�k:Y�٭S��V*;�k�{�,�N�}N�:�@��2���E0��@�P�SRޠ�Z�AV���:eDqZ<'Q8�"���M?���XB��\�|q��m۶Aj9rdnn��sH�iv)���r3 �tt�'	��XȈ�3�}��S%U�L�����IE��\v�$9l4r�
�����q||����k�\[�71�!tf��a�{���i �"��Y�ִF8E��S⫁'`g����4���L.�g�l������X.�庋�֗�̱%{�=.;�s���c��+0��\�9���u�:j�-�	$�#c�i{/�/yY�r�W�K��W�I�y�H�+��gv)�4XA<�&��K���[�2�D�ٿ��J)q�+�J`g�a$����ps��UW]�}��{���K~_j6��ۅB�����i&=g����ք㶘+p�N��L��D��ɺ�y�h)�$bY􍀧b(�!&3����s*��p��H~���:��ږscܶ@ZM?Ts3T�&XSt\���x�����]S�����YPf;��Έe?�m.zk�1Ӭ7y�H4� �Q*��D�3�\��)HY��W���4W�����iΜv��x��8��}���
B��lKt\(��gs5�(A�
w�TRaMQ��(M�������&&&Ɖ����� �U��xJ>�cdb7x/2��C>�,]��E�Ḵ���=(�u�r;�s�����n���)�� z���DYא;u��D��7���D*u#��Q��J9vfZ��l�v��qP_tFX��Zk���J��=�[K�՝�!��1#�J��t.��Mg�Δ��<��0�|I�!�HĿ�i�R%���]���h�E�sB1�:�/���PKe�e��nm�K/�2�KŲ��%Z�2���y��W�/<�AoGrMg�R�k�h$��f��p��|g� ��'��x]LC�IZ��~��<,��i�
%��miq�q`�Q��=�s\$��D��C�(�l��L&9EX���]&��VFT�
fV!�V��� nN�9Bx�D__ށv�c��@���}��׭[�������f�o�s���d��u l��
"z�9��,��)U;�ioo��1f���R+�#-d.�0��0���d�.B`-����^�K�fuz�l�~2���D��;%Ӫ[�,j���ߜ+5��A��e���=� 9��f��`�Eo0Y5;l���'Nlݺ�`tt�W��9���^��W+�#_�@ɽ��Y�̛��]����m����5���'���ܖ�h�/g9���Σ����ߴ���UN���I"jDmT�"�*f3�̄p�a�>{2g����\/�ssnT&]X��{��/�E��K�Q�pa9^Һ�ҧ#e¥Y��w����뤚VN��t�+˶�x��#ٶE��x񊻽>��?�3��}QI�h\������~��b��ӻn]�,WG�^/���^Y}\LCH�1����4�bĖ K��x�wzz��b]�� Y,Į&����}��,�����w�[�	ND��
O�_y�/DŤ4rp�zzz�ؠ �G(5.��43�����H�{jjJ�	��_]6�D��qnv���%������bf��?a�8Mmmm��,U�02^�)���w�\ �w�s&8��	�E�>"��d.����A&	�����%�(��v���d*�J�]�]���_+m~�X��t����m�[��Br7\ݳ�9�qζ��ɬ-�����ϑ�U��\}�K)���U>�,:�tz���1lծY������-ș�������"�Dz��
%vf9=�t��^D��7����痬Q�Yγ ��k,]��g�\vg)�i̥w��S���m!��=��q�]8��d[v����(�M��>Mp�0v�Go�v�T�.��\�K����]b�&[�����`0XV��5RN_�B�=�F�g{�ےrRUBx�h{GG[4����h�'Cָ�ǅ��Egt�>y���� �+g5X����BK�B��p&��&���^�����5@���n���
��� 7a,qC�N�&��#L%��a���5���$c�Wf:�`��+!#`�)&&&���)���.�T,Ց�d�a��ͱ�1�dΛ�t��t�]h�H�ٰ
X/Q�[�����,g���iii���:��xOh�jZ��^������a}9��V���͒Y�رc�ׯ���|%��Ŝ�ș/7��� ��*�KÏ�\���=ې��»T^������*�i���Ԛ�E3�Ǧ�Mo���]��EחD�i����LF�F��X#0�1N�ay력:���?�H��P�"�(�������Er^N��ԋ�'��9��:/JD�.CK��%��	Q�V:�؊�� AS���gCj�U(w���T��	��ۥV�"C���j�MHr�өEƇ��}��"7Tu�JW�Ԃ�%{P��i�0�C+l�����"pC�Q����i�Q�8�c�R6���@ ��ܱ|l9�XqR7z�z��b�aŝ���8�Իg����ax �� �F�y��]D$*�T�wĉs��Yg;�-u�-E�|�hf'e��?ʸa����P틀#c��"�m���9!pu�e�*x����0-��g�`*?��2c��-[�Rc�e3�;L���{������Z���5�����f-�,<s`<W+�ם[Jp�K-�)ä�l$[׈s��Lq�j%'�����Ir��JO�/,:�g��rk.�9djY�'Q�tU�<8Mnv^�|~Y�rȔ�(ۨ|gޙKӨ���J��*9���O�J�NK���+�1�+�Y�P?���l�6ϡsWz��ᖝ�K��8�Q���ns�h@G�kv�db@�՜=�h�x4� �f�8�{-�:[��}�FH�4YS�8R�n�#|1!	1���(�4	/<��(x�D����I�kXن��.ݖ��Ώr��NԭY��M�jO|D���WN�_v�E��#�<�'[A�cGGGYG:-%Y�������9kٶ�j�W�����H��y�`�W�"����
c	��x�]TlzN�~�1x��###�\���8(W*�@����w�z�G�"����۱X)X^�+��ݢ:^�͎��L��c�%�8Vf����U�{-�&K����q�ߏ%Ή��"�[��� [Jؖ����aqҠl��q����{\���-2�BΏ�jrF��wgcU� a�2�(M}�t��?ȗ�+���Re���L�[�cx�b�����ܟ���줐��s�bHc��,�X("�>Ax���؜��t:�4��T�8{8�gE��Z�e���iUNK�<W��߻(S�%Rgo~�,I�T���ys�Ȝ�'%הk����`���=�j��Z�@і���/�4K9��\����;�$�������#���.+��R��hI=6�]LCH/�Sԃ��v�ң��kmm�NAEB���l�/(;?12��!7O�ʾ��Q�{�>.��[��#=n���t�93y~O��|��X�tjj�i�&�7'��H\	(<33�V�,�U���q��\�ƃ�!�w�7�|�3���'�2c}\���ŕ!��8��I'�c�Ȩ_�)Ő��3�J�$�9�kC�şA']��<K ��bX<2lQ�
�ɻ���d��}'���,�����Q�Rd#��ү��-2�����`�s��Fe�v��xr
�|L��`c`gb�r0SqT�ȍ�(/�M\eI	��z���N9=��������<<��$�wRr!;�$���:�Y�A�E�vY޹
2-~����J/8m)�����n�E�?���5�'�Kا�T(�BO\�"�`��\u�$5��E���J��ciOJ��3v��M��R�Ǚ���k�}ۡp�=�:ճ�X��9�����1��DS5��!�p��\#@}xM3�͐�M�)z�PWJ��X�E�Bi���q��E�ǣ�J��LJ`���l�P���O�,n����Cg��of�s����L���L���>�І�҄���*�F��m�x?~|``@��5pk
�-�� ���ǥ���5���Z���f�"����aX�J3�CN�g\��Ӄ�NOO�xS�D���9<"CCNv�3�N��paaAG)M�/F��F�D�g p���H0�D"���8�i��:�}u�Df��GFF����p�n&�lr�?Ù'�4)��*�a�t�--��8�½Syc�8�_���;)�K�íx�I.x��r��!ЕD+��EV�3"$WDF�����"R�b�xX(���^�.�3�,.�\EtF��?�$�Uh�=�)�������P��J�ĳ
�֭[��>,�'�~.�Æ�
@N��_!�N+�w�μj����3$K��VW��)�e��T�"]��&D���u���T��I���Ƌ��h7B-FcغiQ�\��WC1���R~V��N(�g���#@�Q��j�d5PJ����@Ǳ!�,�I�����7�؉�H@t�ղf��!�H�c�JN$r���3��dK���Lv�/���Pkt�t�Wj�^'D�)Q�����S����Tz&��a���t`���r]8R4���,�E�獾J3!��}��J��̞*��6��xp�9Ep��<��R�p�������j�]Wh
 bio�s(�6�_���e���#G�� �����M�	Yv��w*�b|&������Lie{C�Dc���L2�\sWE���!�/����������l1��5���^�%��<i�\�8����\j���k֬a�8��������xX@�S��*6���`�����&En�[���38<��b>C�$}��C���333���|O^#�~��r��B&�S��ن��$Ē��$l�SK�kM�߈��J&�z��]/@U]�^k�Saq5�m���`�H�%�RF`�Ox�A��h2Æ���!}P*�Z0V�/X&\kM�.\�7a>C����#˲�;IA])#���9�!<�����^ڨN��˭���x���k׮Ŗ�y��E��1����\�N{Oz�%I���cq�$�9ʖ3��rv;�������(~kt�mJ	�Iq&��9�d��4k����1e\N��q�C��Q/���$=�4��/��7%}�rz���38���]i������:�I���2N�W�I���f������rRޜ�����R뢏9�g-��cc�]�/\�P��GHE���l��#{<�w�O�e`Q�ᱤ:��ʳ,�Yʅ���k%*�s���7����k��6��X�xU��,cŁ1�'<�I�R�"B�`�D?1�Tv�\���X9�;�\n�$� τ�5�N)i¦V����3s�ԣ�T����xH�-ٖ��"�7�U� �E/�2!�]XE�۔թ��3E�������hdtl�p�م"�Np��n@h )�K�L�.~D���ă��.Бn#C(���b�����T�*]�h����7��Z�T=|����xkoW�Sc���P@R�����N����S��Z��
���J��Y;�`�����FP�T�z��<��O=%�V�8�����'�� �Ö�'���t��A��2�	�/Hq䴬"U�S�$ekz��0D�5uś�<w��<�l?�"\��E��R�����d	p����ģ����da1�*nP3<<�y`���a ����_v�ӈ�f;A5/3�x��s��TD�?n.?{��ٷ��V��ZZZ�����$	�:�C�I,V�W���D�-��q�T$r����mH���"�d��H�ժ��Sm��X*�Ɲ������$ܬPv��}��4��f��eJ���k�)���G#��r�{�q\�5��XqiQH�1@�s/m�QZj��/%EX����o^�Ze��\%��l�qΜ��m	Uq�8����=�0��і����L��`�!�2 �M��)���D0˖Ɲ�ZV=��w$�r��0��)Av�H;y2�ӹ^2�����O~�#��8<N>|�Y ��`�d#Zi�8��V׻�M;i��N�'����Pa���8p��Bl�Hیϔl
�Q�8���[�V�;��z��曷oߎ�k׮��zR��m��U��j8��ĿrIwSn�;:����j�3888>>.�}f��*�,��c-��������6l`:Mv��-Z�O��sϞ�O�?p�CADT�&�ϖ��ӽV�/.=@�����EæUD�(��f�P��D�-ކt�[&�*�8�g/��E�tlc�Y/������;]�p�8m�^1��|�\�C��o/k�^d�8gGU�������jͤ?m5k��뛘=p�����dKtݺu�b��yVzD�Vq�>���ۖ^*A����m-��tƴݭW��Up�X��ˇ�LH�ƺPC^/�~�� c�(K�8���x*&Sh(LV�[U�Q��.��8��vF��4(�K���� ^��/�Y]�����9�N����b����4��t�ȑ#��^����P#�����ā�o`�LNN�5���!�﹙�S��w
X�pRʦ.�UHL�dtt���4�j�u�
����?1EA6�ş�·�����!�>T�2p�괻a�������V�T&p%	���E;���P��B�_0{�<�c}<cܝ���q<���q�ӝ1?ڦM�:;;��/�_�������K_����_|�E,,l��G�b����'O>|xdd���t�o�֙s�\;����i�;�[�c �F� [zQ#Ev�/�s���������^�!���a�-�E�E�:�ڪXGk[k���������PK�{ 	����^��'���@���������{����|���<绎t�K3]�-Q��2�C�ǟr�0�?Y�b��"S�H�N��1����T��q}P�T�(�9��θ�*PιՎ�ز��ҽ���x*WJ����{TDT5�Q��+}k)��
����z�Pn%�+F�@��ЫD�&��c�ZS_k�B�T;TvQԓF�ի�����ک� J#	�~��^�ꦪ_6e_�Ɨ)�v)��iʔ�W��2HiQa�oΞ=��e�ђѦ��aŎ�Bh5]H��������;[�W^�����nl'd�ǫ������
~4����ɹ���G���4�`ZL&KlzC�h�?�����/|����{q��5zyS���K=�ТA�U�]7F�`89ܷ/��J���>\��'�M�>��#��NZ��l�y�mD}q��@B��y}<)�����[O�i��bq�Z�������< c���V�����6+�\���S�g����a�x�>j%-�������bxB65��LQ�T{zZ����.3F=GJ��9+�!h��]��:�[�_
�7�KT������Ș��Z���2�~x<���DqbgF,�� ���M��7�hT�Sh[XJ@���T�\V�3*����@��A�� e�U~m#�B;�>FlJ���&$$ U�yy{��T"��_l�K4�iaD�A��޾��,bfVg�7xGbنR��~BB.XVV�g�$ 9��'��e&CV@��L�2�qiii j���_y���?
���o����1Q�
���{뭷@�T8�
8<�OʕG�����6�OP������1P���vM����*�Q�-@LC@?d����{�=�����,_�\s�JNf�9���#9rOѱcG���3g�����?���
���է'؍B+�"ʓɺ�\���*�y�~�SU�x}�e��6���
<O��n�tfT!�]����zAb1��]�����%��"]����ڵk)���������4��OLW�B�xH�N��~^^�:�QN���B{O���"�P$��KOOǟ�����Μ[U M����veoz����r�X�~��N\\$��!e,��Ar�0�Kߠ�sز��5�<��9��s���XM�A���9!�/2���*P�r��1<)F���#��/�w��d�6bhrRR]}]��m��.�/����/��h�a��]�(����Z���k�!E�3���;�.�-�4'���Y����[ �T<���&)1[X��r�T���@���`vv�N���R�<�.�*11�K1����m'~v1M����vz�Ĕ�Rr�pB܁�j/{->�u(h4�2~��T�=��b'���P ,.>d�ƴ��d�������U�����M�M�r���DHO΀� ���� pYm�8]�F���	c�Dȇ�T�cc�(|�w�s��L����q:]P��y�Y"1�PxRSm8�6���U�X2�.�4�{@�Ḣ}�}�[�;w���Y3�ȉ�VAi���!@�5Rg��h���**a�R��}���.�z {_�=��z�eQ�X�aI�a�!l�I:T
��	C��10o�����N@�BOz8x��:c�ٚ���b0����h�(��Ѥ��ѣ��\V��VT�UUW�C�E�q��XxL0�a����W�N~(��Z�*�*q*F�;��MB�~����W��f�U�;t�O�ݣ�y��ꫯ���]�t���F�����0c��v��믿�d�O��O;%]O^
[���TVV��'el-��bADH��b�Tau ���Be�o�H�[�>a=�
����999������x'))	��U#�oӦg� ���}A����0��ۿ?��AO�\/�%Q;�B1��cHx��������[<M�t�H������F���.�������F�a��pS2�SQ#0�XSN�ZH��%������/�9͏�щ�J)QgD�F�����/��rH��9y����?;b�Ν�B۷o�ꫂ%M�0'�Հ�^.C�0-xv��F���������w��W���T�A�̓A2I�0�yj�⇕�I����a_��'f���a�<��9��S�m�s���P��p���P�T�K��q�F�Cm
$��7vm�����;��}z��ZL~���'�����<�o��������{����>���o;v�&$qÆ����0H�NՓp2z���9^�����x���/�sA1bg�}�II)���:@�D��՗_qe��~om�gܸ0W�SEv����k���ZPj�g˅�پ��:c��bČE5��L�o�>�+�w���;u
�> ���p����0,H�d6 ��-/�n��!0Iqδ����
�#G��.���HTK�@+4�?"D�*�zT+((ؼu{NN�����ܡS��ٝʪj�^������G;�=^gß��!~�g#��Ť�|�˖~���6����r�~��^_XP�h�$&ڜ��p���qc(���[S[#7r�ᰱ�
Φ=��fkp�Ғ��J�]xIMF����,<w4�<�b��J:��,���ת�H�������@�l�4�5m�~<.Ԩ���x�nݺ��ݻWF�9$4Z�6��s��W^y�cF��ﭮ��;k׭^�t��݀Hx�����,B!z�8�F��MV�
���$~��WTr̬ά�5�~ƌ�Ǐ�bUWU9mނ���o�z��#@~`� m+���_L��x�b�;���l׮8�+u�ވ�]�\m�8NA��+=qv�S�g|�|E��O�8�\\|h���BEI-_�b >�[o۶���c��y�#G���b�������&�ʄ�
"��c@aҤI��?��O[�l���6����$Fg��3���,���w}ᦦ��t�)�i���I@�~i�ar��ݪ*]�e���mt�b*���O��+�g��=s�L�\��3~��=����F���ddd\w�u�:u�������������������?��S�4E�[��DX��P� *���=���-eɫ���Q쓪7��ʥ�D2	��"d������n�W�?�)@��\zP�	��g���H�����J�Tsa�����*�*��F���Չi)��
b� �`���bT��>�IA��������D�+���=�m�u�qfS( 2�lW��rl��>�l���_/��*]�&Lx��z��%Y��d2,Z�ɜ9sV�^��!۸���㙉���ٝ��SA�ٳg�֭|(
�Y�b�bI,b��+V��/O>"1	�	�7z�]w��ܳ/�ۿ�j�àH��Ik����R��o# G,���	��i�����I�p�P(+������A��
��O�4�;lס����(��#eŇJJKKa���K�7Nj��{i|?D(���!ܺu���6=�fKn�f`�~�����5��O�`w��{H�U�����Z3�~N�! /c�b�������:�tΨ��+r�����d��`�J�OT�C���	���أ��d�N�C���X�Ғ��[�������n��A��{��+�;�q����Wlٴ�@A�A3�P~�I]_������sY�[�UTN|�ϯ�y#��Ŵ����1�܈����%� ;��Ç3��KB7���۱cǇz��&�G�<Mo�H�w�ܹE��[�J���e���6}��+����믿|��/_�>����ٕ��Q]SM��+ Bi�]1(���5jެ������C��<�.��=GI�!��A���'0hР��S�r��!�b<�qƩZ�0G���Ĵk�:�h�u9�e���C��9ȥTu�(���Fb�[��^��7���o����^@Eg�}6��z��9�9`� �س�:���������芤�����IS��ِ�|O�
�;K�DS0�]�6ڨR\�U�F@J�d���,���kժ{=�Va��;> %�I�۷/�����/�v�i��w߮]��'U}�d�D�O�Kr���������C�>���K�,%��f�?˝6mڭ�ފ�3~��@p�o�����؂�@.3sp#p-na���͛��
:��V�R�d��*���&O�D��"��U�/f��.���M���B�Z�c�����U�_�j�|������^{�������� � D�T�r�2��������O�<��K/���ϟ��Gar�iyq�~f��8)��G��Ā�~�ipW�"��*c�I�t�(e��;`RR��{������رkϞ�S�\�%��w^��ɓ��޽늕˶m�>z�cƌ��Chg֬7f�|�1�*Se:5/ɍ�K��;~�~n�g�(���։vvP�F�8	��!]B��[��}x��#F�	���7�|sBbʟ��SQQ��fu�5����x/ȍvTfQg%���tʎ�����V���Y�N�ٚ��W�h	j�@r4C�aK
$�������A���
�*k� �j��*�*��kԊ�ֳő�߿G�a��\���q��X�
�t�6��Y�v��*1��ȑ���Ԕ$<vu���*A5��Y-�E�|�[-ђC+�*�w��Щcrj�)�RYQ��GLfc8��Ee#�����ގ��_T1Ih�v����4��&��*��d"Z�	j��� ��yEW]=��?|��V�H\I�O��U��K�q<$L�B��d��L��x�/x}LRtB����vYYY� �Q�<9�ޭ�O<q��������F�>�� �P>�翖�����f������ÛS�Nݰa��r� �
�	d��v�N�/1�`#�p|h�P�V�0a=X�C��O��{�����I�M�Ti\���Q-]��w<ǲ��sP�ڵk��kO��kF�����<#�F����6�(lн[�^�za0�7off�4-H���	�օ'��A0���H9(!@c ��¦M�d�����������B/�Y�楗^�My4��
�	���_�}�ݘ�1l�'>��SOᓀ�8�B�|q����	���DB:���*��+��;=v���Ǭ��]tK�N�����֭�5�\s�y�a-X�`ƌ��^}�Փ&M"�Wq��bذa���AE֭[�ϳ����*�f�H��c�@�1K�a'N��r����#��v�m2�6ȊX��X l��O�Q�X���̨6��O�>��%�}`2!�x��w��2��x9u�M��|�=��߅���@��P��C��	3t��
�}��.�%(i�6���Ā�.�D���nYYY��W_�䷢������d&���{@�Ar^y�Hh�Ԙ���l�ܹ34���}P\�-w�bar�^*��|���?3�No.�ڿ??�FLږ-�^}�����S�Lq���m}M|B���C��t���`<�.���S`$K@c۶m۶9���m۶��m��'�~y�3�SS��tݪ.`��h��LzՉ����^�(3|���������G���c�jD�!1��X�fߺ�lf����('5���(��n�?��l��^O�k����~�>��̌g�E��*,���L����δ�����_,��Z�zmu?�:ɂ�B�5�w�R�Ǻ��FS-�0DbXPp������2mM�.�vR,�z��/����dLb��'nl��9{�w|o$�#Gb�u�����%�s�º�E��yhO`����!��?q�(K2IQ��|t�K�6{Q=�j�b���.w���v�˿�sտk۴/(�&0o$�OҐm���ww�\BRk��
T��W$��t��~�	��My�4�u=�e,�WN�	��ڂA�HHd3���u�z���������g�p5��o�wz�ieFoE�+#��x~������k�jd���	���(=�p��v��m�%B1�\M
���,�ͱ"􋎲�5y��f�X��=��z�JO��x�v�98�3�.���?>]�z)����k]������iH������Z�W	���(��d^���f����6^Y�?�rx�~�օ!��NA�d��-s��mګ������^�m騮R���+h��^������l������wM���q�;�*ܵŕ�  �РT0`��_7;Bw��DH�S��4!���	U�4)*BC��j1�5a[�5,�����PB�殻>~;7{C�"�偠�AhhRYh��V�ꭓ"��r���aڔQm X��m�
3�� k>䯡�o��r}1�!gw{�ÚҚX�m^��z�������hH�y�B����|h�W�:A�����Ѣ�IC�5G#�g�UNAb�Jz�qU�pV�F̝�/����;��_��L�h��n?�h������g�V�$�!xN*�IƇd�Dйh�1�@!���E��y�=#Ilb}f!_ON{*cv
���C=���è����C�!\A�PD>�D�B��8|���'�4���<����DR��WT$�u~�3�{�P�FO4a�0����`{���ڊ
(P+##G�ՇLh V�R��X�ʁJ��!�y��0�ذ�����?j4���y���8辟}|�m�y��_�W��>$O����I`ς+��S�2�mђn�@c>X՘q�}Ѣ�8ݣ�t�Fh	KlL�%�K����}�;@���aD#L�A ��Y�M$�?'F�ɦ�#��Е	19��4�5���FGDI����r��b�=_���xw[�2_��ZҎ���^���:�,�z�5:���n�V{��T	�|^���'u�'%L�9�'X'�Ť�S�m�0%�ģM�/���lpj��䫆�ʈM��*.�1w��i?��u[MI�Xe���,��u^�x��7�H���><#�y�[�y}�m	�Z��C�ŇyH��C�X�Ξ:��,�c� ��հS)^kġ��A�g�p��[9�h�{�t
����$��*��Ѭu������ -������o�F����cfx������rJ'�z`����|���Z�k�^Wk�1�����T<����&�Z�rI��U���Wj�aE�п�/�x�'�EA�6�����Ļ����t��R>�1V�!dmY��4��ʊ�\o5}RP����檪%���r�����?�g*vQ>�]��$�����$��Ċ�������s�43�|��)�%����_�Z>%�:Qs�>*�I�|�����/q|�h�!B(���H"i4�����ҋ5}%����n���U�V�} ,a�`/k+������L>����`e �l�/|p����l./o.��x �f���H�-=����o��#���F��ƻS0��Zm0F,��<s�<V��@0��> QJ�<85�1�?��_Q��̛��t�l�X6[a_?����v���Ȁʼ����=N���s�8�Џh5��_��ll��h<p�&�Db��u\
���G �#\L����2O�D�;�3��]| i�9E�>��PZ���
�Ea��F3����ժ �V�ǑP��\�fz�~��Pj��Zas;�IS�Ux]o��p�4�ӑ[h��x� �V�"�±j�M��2��mFr�0�[���0��w�[��+妒o�o
Yy��~/�ֵ�P�ۋ�?^�����p�h�~ 9����#ubC��:}���~q#Rwh8��C���&�h�(ӍѼ-����Ò�������0��t7j6l>���f!��a�EH���"�/l��p��(��߫����Ǘ�ˋ�Ӵ\AWtB~+ĦA@!��l��,&{�F�*���pt��e?:��N:F�Z;<�.Ɲ��UM�6 ���?M�D�u�x����B�_6������#�G��.�QU���ƈ޲?��ؠ�RgE��}�g�>�wi�_!i�� \�X'�0twÃ���,Ѵs�V�������Zlҷ:�cj�/��C�*�2y�AO*`�4٢��V�����W�8�k\ѽ�[��=�>h�)�1W��U+���Ք/V0�Nu6&��ď�f���Q��ʙC�ܼ�Hb�+ءZ-�W�6k��L��P�k�B�E����x)��S�����&�#Ok���q{��ӷJU5��$��q8�H:�@�����/�p�E=�++�R6`@�&w�~2�XY��������l���2\�,r2$^	 D@f!����
я�H��H�2�����t�3�$	ǌJ����Zf��Ւ-ȡ3���z\GA��:�@SC�"�f����{�@�j�5`����z��v���-Mn!D��{�,��	�4n�G�S�nn\�a0���T���}OJ3�γ��p	�=ep,�b� �E�ε���0$�0��Ҳ��$GR�����]��9�*�c���?z\C�4ۣu'͖�ʐl8�[n��qZ�e�$�,C�KRh5	޹3,��(S����� � �vWW���JkH�;����`x#l�y-�T�&sߗ���v�����NZZZX]���ӌ
�|_���\�H���X�d� 8 B�Z��]Pj�J���T�:	,�����[�I%�>�WX1X��zX=xh�6�͸��]�vou��-��7��?�$ږ/7���p`C�����L"���P�Kf���F'��HC�?��o:�ć����Ti6�Q=`�.CZns�\��P��C�BQ�@G3�_e�q�1��4�PZ���=ւ��!Ϟ_�&:>�Ke�	OШ�˶nn�H{~��7ꮰ�R�(����U �~��9�Gm:������F[Si^�|�Je�����$$�E��!X\Bř!�ii{��(t��߆�� ����NP����䤹bX����ݓ\���%mT��>�9}�*�;]NA�9�\P� ����.���IM�?T���~���Ч���A!BȂ��k�j��(�h0r�A����W�-���k����|�xp��cf�it$�2p��{��j�pJ���Pmcx�*�������[1��rj�HG�����+��k���b�Y�޻�bw`=5�s�XI�{q��]�qҙrP��6��(�֋�ؕ��I$����}�"�����XXR��k��F�1E�v�~�~�B�	������vfj8[��?�Q���
> #���*��b��}�X��KJʡ���(/h�h��%.��F0�8<������|�K�į�R��R��ٴ�W}T��x��A����S�`��u؇0��vn>5-mt���N�_�6܄8�3QvW��}l�+��4�^�N�P�r�gr3�����9�XpH�C���&q��T�������BjEmm6���z	Oa�i���S�Lr��.I�l��W,�:u��)�����������v�-e�R'��l�U�#��OIz���Q�S�PJq|���M�ќ�$ĵ��Df�
rN�_�O�������&�ؼ�-�T�����OYR#[4F粴4N���g�VT�(X@���o'����͓�A��t��f *���1æ���������ٸp�
��e�qR��W��Eo��i.�����ӝ���to{1��+��;a�1��L=@������Yb�Z>N���z�'���5�S���"����ƪW�cZ���l�i񶔪�?����6\�A�! h#]B\�M�	|>,�뺑Qt�|����^�t=��8��¼��������EB�C�',�6�S���Q���!�l�r1c��	�Q�EB�蹶uSW",[�t��݀���܎������ x����p1�����[��z%h���D`�'�0Ų|Х�V�		�y3��E0;��[�\�D��],W�2�$��Hƅ7�/����������1�W�LrA�p@7��.~�� A������F���4��ڬJ�<��h��)�v*���"̓��t���=~3��VK.�腓,$��2��`q�족vGX�4���!�����@:2���e/��K�0��*��
5�?���0C3�Y�����"�s;���G���(־법T2@�����r��zĮM|s/��`�f���ZC;��Y^��N�z�����'2OP�u�n8�N𣙋��;�I��t��[�8�b�~ez��q�5E�8�6�<�@ۦ6�2,��H(�d�g��?�<�w?���7����t!�i}�/�?X�:�;���v
".'+��B������_�i �Ux5���րQ���=���Ï�,��Q��$è~Z3��߿J!�xF����<|��kU�8���BCs��O���|����y=�OO\� �|�1���Ɏ8<k����"s����~(��wM�� � ���H��K�wm0v]4��nT���L�<�<�B��'���Ɲ�
$v�S]�TU\��ΈO��t����f�56��ID�LQ��k���{�vx|?FP��T DǾ^�)�}P��Cy+w?Qp�'_�<D�z�|���:e���
Mܤ'��/�%���ㄪ�G��]����&zeCýF3�r���D ��gw���+��$�����X8կy��~��{��;�N:ʮ�-�p�Sl;H<-�%�����ib��i�_���$�-Le�ȼ��7�UA�;��i��)h��,�7�vr�yw`����胷ӁO��JF�#�.�dt2oĩ��	�A�2'I諦y���a���Ѥ���+��6����o�/
%..�0b�͐�S_����r��yꟑ�������}�	Yq����65�'�D9y��>U�Xv���$B��RY�oe�2���.��W9����FN|Y+.�^t�d��֕��^Xխ�u5�&�JN�*�u���Y>�;��è�U���+嚐H07'�}��H��"Z����X,�MA�L��`�М!��^*�T�=�l�rJO����	s�a�t�w?.S^VVk�G�ߨm��X1|c�*5�V�3��~��Kti�b�o�$d��Svu(�I��`C #���{�%;;W�2.U�VY��rָ��1�f�dZ�m��.�5���*�^(�_e�F��4��%��V���T���hf���K-�c���S�MmK"�8/r{!j��M�觢�(ڪ�v�����R|]4���"L�ΆU�g]$����ٮ�ւ�a��8�yj,���uP<�b5�{$;ZZ}��\�~ �{�7�E�pwt.�%Ǡ��L~�����,�1�a�T�}��S�`T@����D@d
��r�3 ��!�Ts'Mۋ>M}\z��������[m���0W|�����Z���x�R�Z"�4�w���qmRZ]� ��Ga����$�zw�Ĵ'�u���t�`m��ϴ�^���#�n��ՔOqpUA��{�6�ʴ��<Z��`�P��@/��z���3o;�`Y�y�O��v�����˱��Y�\�4�b���tx��ye]Ń��t$4���d5���>�,�4�}�/Q��D<�K���o��L_/t��,�u��5�#�wX�ށ�=��x\Ϋm����6�9����s=�I�l�ف�bg�eY���-7����b&�&X�Y���E�.��/�l_�m�pf^�Q6�*�am�xZ+��᛹r�����'��P��}7bCAA��Y>~�Z�]
�)���y@��4���2W'��@���U�mS��BH�Xk�g'��p��0�ż�[>w��-,26���
���!�vNG�0a,�PP_Qon���}�F"NV6a,��/��E�yX� �@ �b͸)����f䫷���z�j��o~_��G���)��,7d,H�g���Ⱦ�����[�􆺧q�_==~���hql�E���
�J\@%((��ƔT��z�ų܈<�:��]������Qr�4��/��V�$%�[��!���ٱ4�5�8SnI��n�L� F��dE�Wa%1�d��da���k��TM�G�B3�j�$���򋡽��
�U��2��gk-�6�v���;Ұ�xq�j�ۥq�����/��?, ���5���:ϛ]a>��6�L}M�\ܹ����EY�����Ϲ���|��3Y��j���e���'A����m#0a�f�|��l2����-	� "-:`2�����v��}|���c�D8�6e?��H1_��E��ޝ�B�Xa��|ȗI����N� ,�I� �X����zBH�b!�;��1�z2z,�/�o���U�����V2�������_����Y�{�	[�a���α-����{�<��ZD*4�������E}:<0KtD�2sit$]� �A�P�-C�(�:�u�t�|�x��u�.������:�E"y�J6Ā��_��zՓ���[��`F�R�LK�2��Or!��Dg/��_5�~����i��r$�Zy���̃w��_n�	^E�ܮ�B_q��80q�|~�K�K{9�X��ϭ��d�V�!���H�Od�A�����&\0���4�6A�������ĬM�h�W�n�d^*H�ٗ�iow��jо��7���OV��8��g&K��mp�?���M?�1.�8���-+��Q)�T2��I�h�b'�A���(R�7
��y��.�C3WRd�>�%����;,)�j\,!�S��a�ќ��vE'P!ˀ�/��b6�;��gx~���7�(hO�s@{!>y���Ymr���<��>�V�U��ӹ��Z�b�����N���3�7��4 T�^ͧ3�}�{�����(mMp��Ft��0����#bs���N������}�h�K5���\d�<�.�%��3m�����ї��`����G��!E[�]�:��Kя���B�-�,�;_�?���������)_�RՄ7R�P��@�,�������|C5w�Tc{�;�|���ŕ[��?�ZlV�x-T���slk�@
L�űk@b��r7�X�YÍd�����uA�m���=k�ߟq/�@
���贚-��㭅�G`&��jf����o�5Xd_�n�.7Eo�f¶}����g�bI�W@�6�8t՞��*�Я8��/b���2ݺ���7�dX�2u��3O 7��DGF�*�#*��`B�5ӱ)(.�<�jۯ��_y�=��HqҠ�G ���,�4��V綇ɏ8V�p
Lטa]/.�h\���T���*J����=�g���JK%�� �(����,:���@A9|�b����p��<����p�uZdo��S��H���V�`�$԰��f��i����?����x��R=_ݺT��<�4t��g�/������kjkk�i�)[�pQ@!�Z�rA8�P�a!�}�_?�:�r��	I�@P4�f=��o���<��A��{M���ʩ��0�gsڍt�yP�O�YVT�V�D[d�t�&�%9>+���9�.�*��bY����|n'�|�|V���<��Q9�������-ĉ2z��@�B2�������t��f�,�.����zRo���h�I��'�6�ЩI9M�X� s�@K��>�'%�Ik��x=T��ǝfZD�̌,R�n���C�����^Rqm*b��̿�>t�z��`��d���jz�y�w����>c2�xW)�OFt�4 _�֮_�t\�M�2�,��q��!�Ӳ!O��u�X2�h(L�ű��)��G��7Z`��7������W#�=��Dg�z��gU���q"��҈G�$��o{ ���|���8C5�Q�6��9'S��V���c�^i��%����A�6*��E5�a<��%pN���em�h����M�Q��#�XYmݰ]\[;4b���`g���~�Ӣ�|��YL�ע���a)����6yJ>�r�L���j0	�q�0��2t@����<��s4�#���Y���}rm���Aw�1Ū1�p�#�-#?�Zl�������&'v�J2b�kH��I/��⾟feFy�0�	�߰/�����"Ug���u���/�tX-غ�[�k�R,�4Vj��0b~��_J1<?��p�����o��̦j�ʅ=9�쑓����,dK�̕�ɰV�h8���a�����������+nN'�I���Ӊi�W�؉V|	
�QG@T�&����n�z�Ҽ���Ry]�d�+gKӝ#��U���A� �YGW�����W�j[J����}V�i'/5ߟj;m�QG,��HIt/A=i�eq�K&W�����{_�z� >��r�f����H�LE[���)D'M��y���!D���Ьe��Fy�v���n���˓):s�&r@�[y��_�~b3�p���������h�YOϥ�>�}a#K��у�`eu���q��u���|���U�n�!�6�0�V���B_��Lu슚��p�H���'�~(�@4x�p��㽊��K�x@]
�7*$T\��x̗����ȯ����?����ArbLLa���&7.W�o=�;n�v;~�5�{����[�K{?�s����pvq�����3:�P99է7hP8�	�:i�2��f�3�3�X��HZ�S�x��?gsSh;VLT"8�_9����*.���㘠&t����/@��1MvG�-q�4]�\��l�<|��%?W~����/�k7a������q�A���G!�{��ֺ��>�����
笥������]TJ��|�&��1*�Z�IG/���o{���!��NVOV�1���,e�C��~(m�����ڡ;� ��l�z���NlO�Z�iOR9L*l%�
(�̝�엥���p쐰�C*N�{JF=����TM,�4��� �W�㪮��v| ���:��Y��C��բ;�j�v�oq�q:f_v4���ft��)ƃg��L��v^1��׃xA�urZO���6ko�@����Tf�JQψ`�ן��ri�B���V���NN�i�)3��m� ��v���W���G��P��<�[�Q�sj�M��Hɏ���v��bE���\h׽[�
��k�5��H��5PBx�-�Q�N�P� @0'�4d�6>�;2����:�\���VBV���1-5��ˁ8�f��_TE��&���Ql����׺������U���p�a��Hb�l����B
�� ᑄe�۬^�7C�q�u U� ��_�r���j8�6�G�iO�xR=uc�
\6��2�X���'(���ѓ譣#�����)���,��|�.�+�I%����9}�=�/��zp鴄f�;�n��yXL9�Q���޸uzf������+WM�A(%�p׹�O�N�4�?�W�.n�$>�7��qOψ���@-7�hI��@��E�)g���Ro?��9[ꁭ��lm�;5�����^��vC��"��2P�s^�i��6FΟ�ƖD�V��H�ʌ����$�B�R����6�
�.��4f6���Lu +�a��zZ�J��Y��~�kk�߰u�	��z^�o���=Zqu
هc!��a~�W��	������9��N@E����vz(�Mc|��0�=c�F�����CXz�eR>��J ��&�7�ۨ�x>S+�;���`I�y�z'Rt�蛻c�$m��l�l�4���5W� �b���G��|�\~~������`V_����m]�n�!.e&���%�K�6n48���b� �[�d����Q\|�~��ר�������;;�Nƈ����q��#���b���^�n��󼧒z� ^���2�~l.�Uբ����񱥈4 �j���q�j��{�4ƹ�h�ƦZ�G�7m�Z�Ru4�/�_�3z�~�HA�*aF��PD����Ȑ��%����~=-Ϸ�^7��|ٮG%��_�|����<fֆs%���x���=�U&�u._?���d�Z�~��۩��c��g��k���;���z��B����p�3"c��98�z��`,��CNyG ��n����m�6��n��@Î)Øc���:dؒ*�~}�	D6���,eTO[[zl�?4��z_vaO3˿��kΔ���(��r(5�Gig���������7F����[������F�d�����������~�)���(�	��أz;�x���%$�(0��i����*�(�+�W'���Xo�[��3��|��ԚH�Y4R]�H�<*b���i���̖V��dL��G�g�y[6�Z&�<w���8)��R��MYK�m�U�����a��	Bc��v�y9�3h��O���$��'�t�"�s���d�*��8�nד��c����:#Ȗd��n��l��Fq�����ov1~$����Yf+b]�j�,Oˍ���/��OM.k��Ȳz�D����k~��<���%d�E�K���R{�Xmu	�1�'�nx �A��~�ESk�5�⼞~{�G��E�2�O��(����q�_�G���1��y�����PL.����p�����;v��<H��E{o����X����¤�[�F�=nG2���+��������%2
Ϟ�}�tFa���Nc�� Ϧ&�k�c
+�����92C�W�8e�Xժt�Z��6[I�"y��)�Z��&&�=���G��%���DT��*J�}��h���z"����lf�͡h����i48�U�qz<[��d����r*�1.�_��s�D��GJtE����fS���{mի F�P�Z�L�� )�K)���]�<g����Z�(g�/�`!U��I���.�	jA��[�������T@}�z�m��1B��2�U�Z t��2U��R*_���y�x�G$�0�u�ިm*0o��������N����.��!D�
a�N��u^wO`�&� OY��
�����ˌ��O8����@�����=�s>Wף�q�S󃛁��C�uhd���g`1]�U ���b�2Q���*�$�B�gLC�KbX�i0rz,�p�Gb���^��f���?����F��n�;sǵ�}]����Y�����Z.�,��D�_�^��ϸ\~C>�a
�ų���W*SfQ��-:.<$^tnr���!�D��>��'��͛�L�s�p�F�v�V�� (�m"��d���a��/�T����@&�C�7e��ŔW�� 5�0I���PC8/��[V��Iw�au��R�
�F��Xܭ��'�ޟF�� Ղ�@eJ��]+EșK�6���HU/ͧ�j��^4ƀ�&P���+�,{;J7V�{��f����؟�����ר2���ei��b�8��q����}3���;��x�/������t���!<��i�K:��o�h�`��hJX_���h��?��ڃ�R��������Y�خr-}��l*M���t"�\�L.0gy��98�T&{�,i��/q,i�j�E �
b�ĝԘ��A����brj
�����^O҉�͂	�H�0���r�b:��x��]K�>�������W��3!&B�a�E�ӓ�%�fh��]^s����^���A�<�w��{i�A�>x�O���� ����b;	�r�	<L�����S�K���6�m���t:���N�����J����V髖�  ����j�Pf�x��չ,ŀn�ib���`��#���*����?��l���7X�O@����%�f �@�;[�����~%܅38�8�%i�4�`Ֆ�k7�������E b���s��Ă!��*B@�3��ƹ{�T �"d�u����kT�J�ڶ�`�6��f��o�����,�E/��$�	 ���z=;����D.�F^��Q��	�{�F<e.N.W��4�a.)����n;7�����c�Ҳ� ���[d�]�b�	��a[��N���`�O\���@Za�7[�>)����~��e�^
�E�h��4���B��p�x;!ʆ=���f$�L��y�*S�1π�[���z�6�1���/��_]]�377��˕233;���w[�U��E�C�ɋ�)A�B�J�,�D&��M�uY�g!e3n���P�J
�[|[ �@-G�ZO�tz��¤!����zۏ�<���|��6^Qjb��񘜢�n��߫�]Qv��Fа!�����,A�A'��ǒU$�<h�C�ë�wEn�/-������.�pُI�Åԅ�	UQ1}����~Z��%}�����
�紘�����h���l�+u}��T6۰�HQW���'�wW��2́lz_s,�8WUL�(����]Sؒr��<:{�@F���g ෺u�]6g����)�v��S��)�f:��u�sZ�_@�N��C޼"��f��ߟ8�����v^۶o�����]�$��'�yt :��k)���r�|{�
��4��`��0ϳc�+*�0�����Z�яH֋;�E����$ZP����UU�1a��;ù K� @��%�<�=�-�X윔]�`&��H���e��&I� E��.ȏ��L+�9NX��Bq��ɔ+��̂ �q���ZgB��ڹ��:E�s����������}g��(��KJ�E>��R�e����l����g�5t�2O'���� t�%#'��ƚX�g�Q��h&�YR�B��f�D ���N��X��D̀��h������̉U�6�(����DWN�Gč%y@a���jnFˈ��X����p����Q.o�h�bI���3X$�J�ߓ�}<`�����t(WB�� ���3�u��Etgg$'��]x\4�1t]4������ݼ��F �E��P��� %�
'L��P����Կ�?]�U;ܴ�X[��17���4�O��V���F�{LgЏ�J6�x=LF���{��b׃�	�>c�{�~[ј4�'�ψ³��|�u��Z$�Q��g0���g~L�w�P��9��t�A:�����O]��tM$<#M1��$�y��4>�L������w�Y���~���9�Fi��a����������4s~��Zj0��A�0�us���+�Ճ7�!5 �`X9�p}�ϳ��X�,�K��];��"O��>�%U�4��d(�9H�U��(�,Ջ����/��	m��� ?��������,�^�~y)�\Ӻ<�"�?�ɔ	n�\�c�p�1��v��n��EȎ���m�(�+�?���~�G,�*'F�[ߙ��_Z���#��L�#��<,)�)Eޠ��f�t�����Z	V�0��M�SY�n��1����.n��g\l�`R���e�=��qd�����M�ȈYY��������V����ס'ޓm6m�
)+BeW�nu������w�Z7}��
#K��^X�dP�x�:y�Wۄ�]*���������-���]@�J��Ȩ��bL��b�)!{Ά%K_!}Sunc}A�/|��;(�-�V���S�M��KEOë������&A��\����Z�z�*"T{:͒l���Ϭ]�����f&�O�� 413q���z���n���~̥w5&�"�_Іd���o�b��gpp�M�9�]5�X�b�$рU�t3�djk�������g���sɭ���7���e/�*$g�"sgA�|�}K����ma�2P�����Ţ]�j�,���~�s��o��v�����~���-�b.ɴՐ�r0&!Ku
P�0:v���;���m�I���{79=	CD#X��y�n	x�P��᎓�rJjHD�Ո�Y6"�?��ݮP&����E�3�j�of	�[3��|A����n�s��SS:��h���L?��B��BX9(P����[3X��4c���3�ܿ�lu
��,���R'��D��N@v�
A@r���xM=5�@�G�������h��G�|�\,m�:���e?$��g�������i1����LI �ϣ��/�j�F�X`Y(%9��X�/2��\�������MTm������n�*d,��/,�#����(�����Ոo�J���v��ę�l�#��G�A22����_�k�ڜFY������O����m�y8<A���p�7������5:�Xb��	:����X�)p��e���O�5 cp��>ȝ�`��o/���.���>F@H�P�b�fdP�����OE��7�j�$G�DR����e��!���`Q`&��u䨤����︵0R֯���>������&d�^^k0ѶŹW�Ҫ�/��*"�[N��m'�%��`��[bL����hy��x	_���E�M1j�&�&�c�!j�;*ޭ�+��?�����t��kԠ���}����ʎ��,��.�3HKHg*� 􊚪��R�����I�W�b��{��q������}�2�O��C�6̭��n�5_��I�����R,G<�K�����s}/0�C�C�йL��+��,�R6ԅى���{�p8<��ޅ������R@A*��BS��g�ߋP�;\����'T9[N�X>8
��� r�5�	~��s�u=a#�T����!��mo��'Hh`=�u�>���=����'$�m�@ގ�稞��gq��+_������fJr������4uH�-��ݥ��d>�2�?����d�VRVfI!�]a2vqx��;�ǂ#���`�xLk�M�7}�t�1��7���k��x=�{
*a���yr�ǷB���ni<ʑ��㘶zz"�1�$<L�F"!|y�/�L �V�c_�b������ͫWքL�hj�����R!	t��Ie�Ç�r�Y6�􊙻m�{a�Tn��@�&���g�R�t�
�}�?��d�ΞC��f�ff��&���.j2|j����@U�8���\�tM�PwɊ��(+3��܀o��A��<e����:YGQ��L8ȸ�JFǉY)'FR��02�EFC�[?лz���rcԫ�r~lQU�mAѦ.�����},C{���TU]��[C�b��j)��� ����@,:������=c~0�j���f$�Q^SCR%n�!��!��l�A�%�+�y�����'����d� X�c:>/��1bk�F=����e�<���h&�_ 4Z�V���IL�E��$siv<����w;��y+b�
�&��"� TK0�]�2y��XЂ�UN��T���u=�/"C-������k���2}Ώ��pY��m}u�Z#��䙀|n��㹹�+�-�?f���Uտ�[l0դ��e�j�?��og���G(A�#׌,�NI~�	ד"�Bf�E�qϚE;���z߻�&���D��=��-��G#���V�-M�*#+����E�fB��np�!z,��4�hS�������'����]����!�OOss��a�� }�RrrrC���a�m�"���ɇ/���4A�����9��q�nn@a�'tt��K �ι�iļt�����S�"�BAa§�P�=����6��q�%�GO"�EΤ���9�{9}R�E)M�����T��~"f�5I���p5G�A�&dW3	�.���s�I����ޛd8�������FK����&����O}cd�)H�z z�;TBVt4db��VA�T���I����Q��0�,Y�Y�'!T�*��w7�����Q/��0�G,�a���\O�﷽�����}Ssy\7���"OQ���U��'�L��F�`��2��`�<�����c$��9����o�r�qe�?��s;�
���viL�A	���)���p
2�ə��a���P'����<o�VPEYYvl���+���^_��PC�ۛ݁�3����D0�7S��+�����xv;V���Žq?MⷜOXL"�u�M�$hd����/sė�6g���i%zй�&B,�NI}C�I\)�E�)�?�α1�f	±���ƶm۶m۶m۶mۼ������g�t�#Ǖޥ��E��ʇ��[�Ն˾�Dr�j�3)�����|��޽����A`�P�=tә�0s9��T^-����au�}�$m�2��3��y�(.��Y�n�\k�L#3b2���`�Ng��z9��/�� �Y�;�ܞzD� �՚ND�.i�niey�@S���$�kkk�i�x
1IYh��Y�~���:���D�� �����;H���<�hzX� ��jic�����l�Uڭ���R����@IC�60<��C3�w9~����G�΁� i�ڞ�ѽ�_<2�E�q��I�o�MK�p)VLe/	y�!`ӷ[$�,���uvj�rldF�F��V�r���}�2&ZkKShz���M����Uu=��Tux��m8?u�RJwn�6����raY�\q�?�.�pP�!�ص[�=<3�qj�{����S3�<�������=>- G���s2���C\��Щ��uy��:W�\3���X`�F����f#\",��_�C=�xR�O�Wt<�y}s�Q��`��iK��(�4/�e��܏���Sf�� �\�?��q;�����x+;���0����8EH��K��g�֖t�>��_���ʪ�x��6D�j��)ty�s�զ���0�����
 ���%ɸ088�P4;Zt���U,k�u~	d+��o��<�0q���A(D�K3���j�UM�H\ �>tbt����r�pKEGa��#qň�uq|\��U�8 ���[��
�6X�i��>��0��T&�ĈmY@�hN_��v�=��Ki?��yQ�LoR
fw�v�vo@Y��6�J�e�We��Q�R~����U�D�Ȯ���\��$�����H�[Sv	�$	ґ$.�by�~o6E��28��h��q����R<�$]�/�X����E��))���n[��o�T�LnR�=�9Pa�����}mwy�٣e?�ݱ��Yp(�ݭR@� |��(ɰ��#�ef�4eV��|�Lpfg"�J[�J���;���0�!�� 7��>�ڦ�J���]������r�(�`�B"�1��$�EW|3�D�I�,*_�5�﷓:�\�}����P+�L0� ����~hZ�_X���ͅ$���Y�T'*�防�� /+�XVMT�Q	1�����pU�%ڮ[�Dϫ�CCsN�2^�Vt3y=`(��U�.V��'�4ؠZ�`3�Q5*��t�zMs�Q;�6�qf�>������A��%'��[Y�ۂ�:/�'�]�ڝ�fI���d����kBa�E;�%I���j�K�n�>��[.7���i���ګ��z���`�e��}>�ν�#9��>�Ɖ��A��ӨTb6���=O�<[cQQ�z7Zn~>���� ��~T$��n��f���!MA7�����t��hA�� ��%a@���(��*�O��@!(.���+M�wNI1a1A{��
>��q!���35\��= u2�'x�q�9�IM6c�J*ԥ��ƭ̻���ZE�D��s?>�@1w_��=c�ny�x��1;�P��3�-�i�{���ёq�yllLߕʌ`�m��������(A�Le�����+oc&B���5���_���u��MBTK`$zM����<J������2iJ�(�T-����"I�G0'�p��������i�&�A���-[�j��F�P�-u\���Q���].��W�M�8F����x��fs�yM'U|�U�(�#�eD��S��M���}��0�5D�p	���D -�v>LKJH܁����Lm}܍��|\w�4
P||���J*O�aϛ��4.���_Tg0x����,L7
 ������ �@)��y��[���h���{�����C��g٨���x&>�E�$w���F�#<S�޵$'�;�������?��t����a�	�U����C�w�����	Zs�A}-������D$����pޟi�+�� ��w�T�������rN~D�ꋉ޹t�@K�Q���Qg��gA�	��n}	g���-Qw��EJ6�(���1��O���	z���1�9~M(�XO�^�9�*�HhK���+�>��`���в>�_�M�O�n6��x
�
4�����<��2�ܫ�@��1xD�H���qt`� 3�䫨$W 'h{����*Knr��_�Ἂb������x|<[ 7�Ҳr��_3͙{�V�phГP&������
r9&/�%'��������;��w6�H����/�F�����p���:S����3R>�Y�0Z_ԭ3�"�5��ѓ;jt�5p�HH����Z(�A�<>��g���3��s"[G<`xyRf�ȁ�|�-XR5�4�{�E���J��ҁ����;?���kܐ>z0(�ޗ���<
���C ����N��&�;��������;��B����d�D"�]�B�(��yL�a�]��aȅ+ �x���S)�fO�N�jP���	D���y����x�[��Lͧ�l��zZ��J7��"���]W�xQ�{�/@S�^�c�
Y�si�͘�T��B\�[-� �,2/�h��,�?��/�Q�1�Vߦψn�d<`0ޟ�30����|z8�?��\LLm��}�\���8������FeŽ�(ŜM�dv�|9��oo��J�؞�l\��SP�A��l�T����Սӌ�Ha3�H��"���D]�=R���)Y�jwu��d�l��B���r`�ȧJ���zh�?-TK��7h�h��?��X;�h��_^6� �0Uz?L�Kmq�	�kLtm�;��K�@ླྀ�ffvn
k��0j2�P�*�Z��p2���j�I�h�ެ�I����:�3?->^��f6�T~)��a�-�W��X�5\�7׬Xڷ|J��˿+j�u����1��|=�ey��0��M�d�)�?L�?��a�/�?��n��G�q"�&(V)��o����)�y9�\�jCYo��kb�}/͔��`$i�,I��{����q{�M�ְ�Cf,���ϗ*Tiu����9�* �)*(��&Q4t|�����q�7�yb�zvlX�'5�+�#��F�X��9�,�)����Ct��)g��zɮ6Z����\b^��0}�Q�cy/@6`�z�����?�G��xh��xLZ�"`Xøa���ЊL.��+�9�Z���8�?*������� 뽣V����.h9�a�����!/-�`L0� ���"\�*��T:ְ�b!׳�C�*Rڥ����K	�����fꊶh�t��H�D�Yy̓~I�?#۞ ��Y+�ۏiW���*�]����p�F���b!F��o�E?�j�Dұ@��>nG ���{�V�W\u,lx�<l1:>5ƫ�3����'�60�l�^����\��<!��w0i�� dY�Xe�
]����5�&���6��c?t�(
�X,��� ��,��1΍�J����L1
�Y>`�:?�m��K���c�\~z�$�Z� Cʕ���v��@�qD���t�?Qӊ����O����Vwl�{ȓ�P��q.)�,탖y!�5xG����C[{+�� ��`"�c�E������'d-@W��1�V�@$���y�����$�7����(kHp����z�o���ot��~��B�`��v����IB���#E[_�=��,&X�:^���tܖ�U�#���F�`%��A�	��9�����k�#���pQ����<L��5����w��F��΍ܫ9�o^/j`�m�P�h�_ź��=Y4�bp>u�G����ɢ7"�K��Pk�x=� g���z��F
��oe�Zy�N�>*AC�/���sL����cOH']���[�*Ӧ���D�M�N��<:,���Ҙ�%�]���Au!�f���;�W���w�'/���'�I=�VM2VA�F9G���,���k	�fo�7V�����q-�K6�6����/5��W�ڢg�tŀ�`�at��yيl%d�R)ŞS�V/DH� ��eF�W�	w�802���������=|L��U_X�؊$1B{?���='�
���&&D�����?���|>/�4���'Ű�К�yͮŏ<�pQg
�{�J�\4����]o�v;3r����z����U҉���ə ���l���U֦�x��e��\Q�x�����w5���dj�����(����+s�fEu��I�@�N�����:7"���1�qɁ��4�������{��â�$�Q�p�ǃ�.�]�U�қ�*�e��'zp�8��p��z���)^�OT����8���&L5�˙Zǟ�ʱ�\/�\����5q=\l��.'O�%P0��A���8��$]5�Z_��S�s�dHb:!M����TD���'��V8-Ņ�J�E�ڈ#�q�E�����x����R��d�p\�:^H�T<�婟RAVc���a�����"�����Ѵ�-RiYƘ���Q��P®�</��	p���� N��-�q>󠮤F����b����zX���i5t��܈KE9R����&�׷[�K�QR-����Tyx����(!VT{�py��[{�ҋ�ۇ��eۗ�0`ZD�\\�T��%{}}�P�˻�)�ZCD�C���\jc!GA��I��v���ҕ.h���AW��@h���O���22J��jw0\���D#��(K����N^@"�B���dWVG:�5���N�F�=��w�g^�dȹW`oW��0�a���o="DЦT&���'���}�UjPeJ��d��צ��ә�﷿���K�s�x܏���*�q�3V$JZ�s����{��Z�m�^��A���!��A�}09���>�1h:N�X��2J�@����6&k<=�tQ\1��F��6�m���ٞ�:=>��m����t4�^nS��i5$�\M3l��B����'�ijf`aa��2``�¶��~�;+A+bEo���C�~�l@��L�A����t7�X,_���Pl�#֕R
�85��vxGZ����<���J�'��I�������L�E)Rɷ3Y�p]hv�~g�"��=�S�ٱ����V ?�,
�M��;�=h]������&����#�9��[���H�n��)
�qy `���V�8���`�\�B� �W���o?���>+��͸ԟ���t5 �K��ʕ�L�$r4Sv�� ߬��۟lr��:�0�&�W`Bt?�b�r?J��-�TsN-�8޶���=[(ٟ���Gʄ>�ydF�8�P�6<T��* M4_�,M�v���7(��
��l�Zc�5b(�*��\iK@����������G�SFI �ױ�n�W
*��7��Qt657��8��>�����k�َ+/ki�8��	�B{�� ̦ݟP=�g��u\�C�5OQTFy�Bz�l�f��l�����0ǎ�<h���|4~d�m�v�,}���
f�\|��Yg2�Y-��|��hͮn9fUm"���i��aL�O��g��xl�fCi���0�%� �,�Ay�!b�@]�s�ٗ��C��2fC����v<��FbG��k47�W�`8:���jy|#�ND'����t����ö�g�����ַ�på�ec��d�f�SI�x��$�_,� R�\-QV�^}��/ײ�>$#�΃��_xWSG6:��u<����o;W�eyu�!������"$�]�)��.��YHM�̒��Z߳����@�� ����BD��
:b��]���2Œ��ǅ��*�ϻ3����f^ +ʫJL��4`OF��b�0�0�7��'f�e)tH*��(S�\�눡���vi�V�n٥v0~k4�_g��i�q��rǧ��I�ʋ�v@����Zx�4_��h�*�ÖN���C�T��S�=���]0cL�M{ל���U0�j�!8�e�i��ׇ����QJ��b	� ��0nd�HIZ�c�U?o �w�p������z����8���U�MϏ��"Rt�,�km+r2���j��׍-���u����CT����m�R`w��]�N�Խ>[��<eD
Uy)Y���|�dh�������h�ӝ� et?��D�&4��G��S]�M���<kL�����8�$ܫz���gu�RPs2����L���>0��&N��DJ�N��J���͝�φԉh��Mi�%�_Fgw�#�Q�?��� ���:f�� �a��D�?����8O���j��Ҋ�m���j�gFy1��L��m�(%.Zi�OwG�)N^`Y7�X���x�3f"G��go�3ٿ2��Lp8;*;�tQ�l��l����_>-��%@����m��(��eHQ�$�es|~!P�e�8�rc~S�J�rн^����s�i���IL���J��9��������}�����_I�i��R�$ϳ���[L�o�dڐ���+�\ w��� ����!N(߷n��TC���5",�7y'�<d r���^4� tR@$ ĩ}(��6����GN���!�����4�΄��	QD����8�PU8|�e�D�M�۳����0���w�Q�-Ȳ=�g�A�
<*+��x^5�m�����VuCU��bz�WL��nĞ3����oga���K=I	�J@����a���V�?��_��W�1!�c�4v��F%�� `��0N��!G�-9�þ��j�M�� �a������v�
�S6�?�gو瞪��Os=Hyݣ����P�~:��8Y�D$8����ٌp.�K�W+H;%�|�����@�������}ް���Y�L��i��Xu�s�i*L�S��	'��������e���J���O(X0l���a`o�4�=�J�����ϞLtE����l�:�E"����~� ��d�t��(��0���D��D��4�������6ʹZ��6KCH�j��\�ĭj9����;�3!���bweV� <a�`�H���`j�//<�m�ϧJ7[��o9?=X���T���g��-!��x�`��#��	1��JC0��x�W~�J���
Z����Җ+�3��-#K�'�^o�6�(('�����U�4ط���{n/��ҩ�gf��u�����*��c��~~�Rb��d�؊�Z��/���m{���?S����� �:|��eSj�۝�N����hCG�'Rh˪�()����j��W�<Øf��H��X��>S����F�߁���G������C1�L�PUl����y?��y�x�`�����M}eG��Ip�4���p�9^���z�����P���PДe�g��c���P)))PQ���HF��r��9�ӁO�'0v*,0"���w�����4V�P���N���"���y�&0ן��x\��:^`�vR�	�2d=|$։����f:�p�c�w�	��E�^H�tm.�>�=���4�����F~�K���9��lu�r��9�"�{R-���&t*������(c��2,�ߵ����Q�4��P�æ����s�8���r|�.3���q�0�u�EK˷������jrX������sޑ�G��.`K��yYn��H4�Q�ݫ;�k���j�Qݰ�yEA��?�Y�U�PL�d�`$O��� *�}�2 j�C;W�n��a�	>/�.�t_�y;/?�������[U�sZz%���2e����Z������J�U�-�Η��i��uqT˲�H��(۰�+??G������lsl)�h	��hl��EU˫��ϥq�4��y�d|SH����h"���i�F�op8��2a���\x2SX�i5o�@�Tx�t��ˏM����~���� ,Q �W�|���������� ��jJH�&1k���f�������NS
��%+A�&w/���k������/fC���~���|��S�R��{y}ލ�t����51�!l�9 I@<l���.�_S�{���s5���T�M��S Kg�ڵ�Fn#8�~�3�|����mS�.0L�1�>2��0����}>�x�BQ�{������Z=u�W�{}��^�r�&�=��8�9p�<�+���"�]m�Q��eJ#z�Oµ��9}7��5_��W��ۧ�s����h�NJ�sD���s&���N؁q/I���].T��E�k*s�+�mp|V�cec�����R� �s�|y̜����+� �����q�Qq�rN5M�������z��WB�Xϛ+�'�Ӟ��b�L�Ջ�F�Д}<�~'��>��.%6.=C����Z�ź�gXk>�ɞXjv�y&~���J[oPI�R�>��?$R�j��W:�����:K*l��ˡ/ �R�z���H��e^�����SNT�{~�"q����VRrdA�{gn��i�@��0Y9i>הN��Â%#\JK�Hy���|[?�=l̸n����O�*�>`M���-m��yrФ�E{�q���ɐ�.B'}�j������d]G�hn���Z�g7;7���Mg���� �ۘ$�Dh��x`|��r�/��l(��`Tm.>~�~|N����~�bYZ���+���+��*���#Ѹ[Kk�s������rW1T`�$��Uv���\u%޸��xE�p89x>O�-������1���9[��x��z>�l�xh�������Ŗ��Ξ�M9	�=��+�cԑ����&�yW�b4��QH��r<��çP�V�����}w�2��%�g�쪬�T嵜h}lE����}=-#�cfn��a��n]<���j�0U�_�	7���d��	رZ������[UI�nƖR�6�\.I��H\3� �>Y���.=I͈3�W^X�� �ef}�w��ˬ��N�P��v�Y2�{z��$N(՝��.U3��/'5��`\B���o�\����O5����aj����ʽ*�������Ῥ4�x�ϛ����c��������:7���;Y'��=}Y����B��'�_�pzR�H���F|D�l���h���N�~L�^V*�Yk��z������ڳ�i^0�h\�潕�L�g��z�H��mCI�l���~��j(������E�B#<4Z�D����"�b�Y��Q>>��\GOAl���o@�O;���N���"I�����s���	A$+�o^�0q��뙬���#�RgN"�\.<�"��6�j���4�_G�H��J$����cq�ô'lN[e_)�+��t���]ց>�9�lbM�E�����S�`m"�b����Ю��g���)j��������1	y[-���25�%b�pr{8i�#B5�:]�T8-&�Lr聵 ���Q���Ng1<��$v��'Ӝ�h �Ƴ+x߷����)����?_/H�{�zT�g���t�
�R�������������������w06����q�����g���3��7U��>�i��Q3��%@Ϭ��C�����/�!y�	Ӣ>�hQ!�2�0>��\��M��K�	�!?�g���U-UӠ�%�d�^@��#!�p]�z%�;:��7SK�*��ف�d�JJ�;�R�|�?Y�̭l��kw�r�x���l�����C�zHJ:�1�31�9�����>�9��1��L�ޚD|�&Se��-�?m��y�EO~[��#Wzp�	I�l�b.Bpdx�� ,������!4��}��^=�^>���5+(ӻ���]�9�L\*��|4�Az�\N`�Ga���_c��v�sg��ݭ�����(Cw��΂��A�̪U:��NA9�ԗ U�C�(�T#Zw*���fR>];=k��(j���ir�@����Lfq����jԇ�
�Ƹ�]J��ϙeB&���ƶ8�@FQ�1��Mr��	�����H�~W]�w�$��`Ĕ���|f��r,-ek��J�k��Pg��)���Jnp��!�L"��"�1�/="�C�O��<	�^�>c�'��gg;�̋�(*z��,�h��5���h0X�W��WO�7ޛ�����`p�<����e�Ʃ|ZPr�"#ԫ�tn��I�<���-^����x*�N��&�H0$��M�ә/r~}^ǵ����9�b^,m��ɬ�� ��\NC�TL��HqxD�W����<��]����ٟ�l����p�,���q~�񉍥(�UPf���o9 *�s�Kd��0%�u\@��A�Z��
9umb�ܝ`4o{��(�"��YX�E(�#B�M^��O'�^Vl�b�r7��Ӥ�@�\���un�N'���Bc��۪�sߧ%�@\,�QND�K+������;������ ��S�#g �#�L���:�8������^=������n�-vӬ��P�O@}v�0�0��:��ha��3)L�Q��-�+�3����OW�
ӿ��s�op�4�v����.Kʪ��C(���mT�9xj<��/�V�{�(��ƕgR4/����z��5_�Wͺ?���+Wc��-d��'�X�y�J��]U����F�mV�W�̬�<_��3�?@f�ģt���DK>�8�`KY>�g��/���l��ž�O��	ٱ�A����D�/E�g^by�"%d��Ku��׶���X{n+���eҘ�>�1�R ��j���=�Ѽo�%i�kȆ{��:zZ�J�,�y�/���>q_j�oǩ�T���\��x�y���{�A��*�4-rH�~�''	+,���5�á����8�v���}!��/1�����&V�~���]�VUE�a��@Z�5l�o�ځ��V��|+"P�m7>@���W���uӞP$R�� �N���[} �K�v�q���=�!B�h������v�ObING�:1�p׊�!(����Tx^�'Q"�58o��� � � ���4[c�IxP�U�8O�����b�ŷ��0�L�D���������~�V_����΀C�����������8B�_M�o?�v��+0s�a� q�G!�����h�r�7r�O2�)k:�a8� �N������1׎�ˑGS�zq��������%�i�F�j~�@H�w�9�/>�����I�d�������PUƌ�-s�ѱ`�c}�A������R�cI�w�L�a��い���d�V��~oL3���O]F���k0�jw�P�Y�7�j�G�x�ko����j\���3�ʊ�u��ju0�-�&\�z��sKKG"��JO������#�\߯���e���I�n���I���lV�{G�k0%������=8��쳛��G �{R�灩���i�c��.������Q�EZ#���\+�����I�Y���*���=r�C-T��`/�Ӓ�/�jI�l�zK�Z��9��}����@�c��$�MihD�����~k�7�k����d���t�apӳB�~Il��;}:�D�\^��1Ows�����g�D��TS��� ��{���ue�=��k��Dv&IuXx��)����lfry��D	���.qw���K�)M��"q�#N�Apy��eſ�lp�^��|�ߧ
���*U]��~p�T����ئ�b*��e�x�B3�� O��R��b��0��{7�����F(��h�)<D�����l��W�;�-^$���ɷ�0/��[tO�����1yG\T��d�{�細��%]E}������m�;#%�@��2A�R�(�������W/���D�//?�1J����St\�~�5	Nv޸��u'S���FK܀�XW�#g�@B�U�ű,���@�ĳ�ֳ�����s�AD�8>OϬ?(M�	��ZH����"�J������r�)�K&�3nt2��?�vF���(�]B"���4�*c�J�q��Jhb;�#��o�tS���y�ذc3dc����t�����X���sR�B��~�� z��d5�� |���q4�}>SQ"\r��h��k�>m�����V��@��`UE4ði(��(��H�>lNA�_�%e\�����%cgSE�x&�m�L��g�I��1Avּ$�*����;��*���2o�v�I�`�M�s7���1]@�Y�iӢ��BI����h=>#k��v�~���n���Y7�6�V)ʬ˻���v����zaa����1�1!�E���SG��Kɒ����Ų�d�|��G����ZO�ݕ	{�h��;^��R��fbD��2ډ� (�j�+|��m�=o=���7������P��@\Ԇ�GW��U����m��5�s�/�]_����3Lґ����F]�ʔ�8��c����V���e�b$�!����3a���Y�t��Z����5|��c\�[+�&�q JwAu"�s�8L�=]�c�� c3��,Q��\�2:���s�3�e���ݯ۾?_��z�F��J6�n� Ӝ7�6�e���ܐ�l��TN��=7�f؄���2
k�f���D
�2y0Q_Z>�*SF��X�ĚԷ�Ar����7�x�P������!���?�F
6֚��a�]���8�k��)H1�r�ƥU�=(ʽ;Uh!O�����D� 35^���l+�"���~+���O��g�3�g����Ф/H9C	#γ�O$_��?��߽�m<S�EY�T����`�
Ƨg(�XH�5�v'15T7�H@����ېB����n�Iv�����]�V�y�q��� b	Kx�H�H��K�@�%D4�	
aa��r�Y9Z^]��)(�SWI� �\��O��j���ݕ�#����$cl�1F�����e.�~�\7��� o!����Sװ���1B@�������_??_��F�޾~p�b��:���t����2L"�MX���i<�b��p&1*ndh����L,&�el��U*��(L����TUP��R�>�5\_�٥����տ0��n>�|Q�s/Y�z�-�{�����yS��p������]j_ ��,�������Y[0���$zL���-%�F�C��>�*%���-LY���`=�8~��]�Q�E�B���� ˗�51�)���-�v�2<���Z^?�o��B���+Ұ�]��ϗ��ܿv�l��/WR&�{�������_U����}��$QP�,w���k/?6\��D�O �u��󢊷����B�
?e]�;ֺq,�j���O��'�.E���!�e,��A�pĳU�\�����ծ����o;����m��ޅ߳��Wc'���o5L�ڌe���.D��@�Ϙi:0]��Y*(��L��cZa�.�_�r@����.%��:�j��f�s���A�N�h~B�7猂�z�,�Q��mGIUՄھ2D��D�nYQ����w�����K��K��+)'��E�f!�M���n�]���n�Ǜ��6J��PMY�߰����e0T^�g�Y��8}<\b@[��a�z۝7�߈ϸdU�G��}h)#��+��
��ظ�ۭ�zl>X���֝��M�h���?�,5��]�Ŋ���Ŏ���'i\�_���/�ﭚE�N>^��Ծ'�4�*��p=���� ��ڣ��6,�zD9(셅��g�̅+F|r�B U	-YO]y&6���8J��6}ʯ��/��.ا(�ӫ-s���5�oo� ��1G@�&�il�9��=ߣ%aC�����w����g�;kϐ��}y?��-6TW�[0 ���n/P�_�Y�����q.v���f����o':�x���.�ݗ��pcF���UC[��Y���3��.����}]~m���7�\���X�G��-$܈]��=)�I�<e����
Z���b�nu.\wv�+	
'�[���so��fhYBG�����o��q�t®i��F(�\��r�L�1�;|������E�ʎ@0��U��6A�!����S�Z��/Ƕ C*��Ȝ��F��*�|5���l�/���5o��|���Ii%�V��gT*��x�6ln�鼦Mh
,�tH��������<(�˧vz})lp�{����i����=�<9�#�(;�v�v�;���f�T 􉶓성p���v ��gS�޽�����202VGvd��ϳ�1�.����()�{���Y/��>Pc���s;g,o��l�R.3�Q=��X�<q��C�=^�$P�r��>��2��.��x�8=z�
ҿ��[;P�@ۀ�ؿ���	��A�-�PJY��"Q�R)��g))�և��2�7A��vK�R!�f]��}�P��?��ĝ)sz����]6�#�2q�
@�f�|��9e�;qK��X6^��''q�6fŶΪ�_���2�he��`<Q\90}�u�uΌW�֥��~9
�;���>0�1W���6d7��Ļ��.�Q�~^._ 2�q�:�@j��i>���G;nE���ؙ�T���64�T.2�xJ���["�ҹ�����!�m�G��ƿ�H�� 2F
��Ak�v��+���Na�
��6�=<��[�D�ֽ��FO@k*��ƛM�S$u}_�>��FJds���d��2!��M� ����:[��XX�YuW�@���.��q�p��7�mu�,~������TF�Hy
���V1/�L�
� ?� y	����Ȝq`�W�\���9#;/�_��d��8y��T�|�|<�Dr����7��m�G�:��#m��1������� �DT'��L��7�ˌЩ� �BJ*��0���ts9Y-N���CΏטA�?,Lq?��#�6i����Ӓ��7�v��ߟ��K-�9eyu���'|��]�؊�?�q��)(Ycr����(svw���=����H�KG�Mp��f��J�r����ן�D��0dOn��������l֔���*f{�K�|-~ �'��@��#���S�8���i-�kkg�k"�����RN��_7����I�&���D��D뛪ɍ�0/`H��媱eFñ�:I#^s�鄥'�S�s���Ƽ�O�~*Z{շ�7�q$E�.���K��Q�A,��ShJ�9S�	`���P0D����M ��X5�)�<��+"G	Ӌ�
���kAy�#�������Q���u���ˤU�,K�5�Lgu��	p� �5���d!N��A|����M@�.��B�5[o�{��v�?8�·�oV�UPX Z�����'�G�j"�3~[j@򮻽������q h�^"��\�� Ʊ��TP��t��&f��L6������F�ɚ��L����yp��w�*y�L'��<д� �D���fX�!\G�J��l�`�p&O�6�у�g�%�a�h�/a��xբ�s��=�$�K*�*A�  O����N*�ᨦX�)�Q!7��{ĉ��֜�$�Dj(!Zc�io옑J��ӧ#�AB%Ƭ�Þ��1��jq��ֈ�����9�z2����e�/vmz��`Cl���e��-W�$�n�r��T�ψa"0вDcX����C8Y���U糆z���|���-���ⵒ��wZ�
>�@����;��᥋&�=.�H���u��F��p����P4�yo{e���
sy���sxِ�X�ω^m�E��в7ڋ�+��&JK���N�5|m��<��C������8�aB:��$�gRÿgy�L�|���I'+���!_@Tm	Q� (���Sjv�s�����������{ ����>��B�����˷��^� �;!9���!!!y �E��L���m7���-�X"��Z8���<���д��Z�	8�-����jP7�E�Υ�>;�I��tV)�|2>?n���u���x�/��c�� ����$
���Q��bm�����E���W�'���a�a��"l�2�4r��]�ڊ���~�-�ZS^�_YNA���㮅�GLr���.��@+ʥH�#���*=���Y!`��w�Ύ��;;�ʞ���2���('�~R�0�w���xxE'#�w�����p4.�D�ׇA�����r�D1�M�^\�*�2V��Oz��J�z��u8JE½��ݑ ��c"uF�ʐB����`�sϥ�M�����r+<��s�����p�<mϽ�I�ý90��j������r���W��rT������g�1��'�������	�53�}���ç�涺�*>`�a�����N,�Z@�q9��]�E~rE�E��s��)g�<4,k'9��|�x�w���z�U���(R��\%0j���ޜh��#�a��Q���o�7$H���?5Wh��ʬ(CD�����>�e�^ܷ�G��4���?ds܏�Gf2����;�
���֓�	P�5:&kbd����$�[&[��^X�܌s�`J+)����c�Zo������˫�� ��B˲�/��`��H����+`+��V���y�YѤ�uB���u�P���L�@G�����%�*�������-�>�'�ⅈ�[[���7�P�Q��2+���.'���ٵ(n]b��5��Lc�o����J<Rъ�$7�SK�H"�`sJ���� t@��|��Ǐ>�X:%� ��������w��[o�3u�+c�L��4D���l����m:#HWU2
���0e�ҙ! ���~��]�p)5iE[��?,�؍�~Ĉg�u	:���%��h�2.�dDΔ!gȜ�����W��i�,,����� �Xx7�X3�g�I�9��X�se�m�,0��	��-Z4x�ಲ2*�C,���?_�Q��D
��E�*0��<�C
;�dW[�Mm�
��e$�7�T��Ì#�#������ڀ��`K9��_|�E:T"�L�$!�XR>o`��ɥ%��,����޽�р����	q�� z�Ѓ��:0�6p��+M�-�?�J�����+3��-qrb���C0�4�����=�vx	9t�XN"D`�y��t*+>]Ím6�m�pmߵ[8m ����$�N��
�H|�T"��' Ƚ_4��(c�W�T(��n����6�� ��uˇ�[�lܴ~���X�X�.%j�̺���._�{xCxx[̀��p	:d��W_Ǩ��Z\�T;&<��#�C�n��ͦ���U��[־
wik���X���bw���Mr��m��j�U W����̿_p����J�
�E3��ԭ{�Ce�� ���Ʌ3�W�,/���[+�����O	���W��m�jU�����[��M���a�����;񤓔���P���?�,EA�d2�|V{MQZ���=W��y��>�0��!8�0ݶZrI�6�~�/��-x���WO�:�_�⩧�<pP]Uuyyiq�Z���;v��5�o?fNgk<Ҿ6�
x}�e�^ӝM��Ca�"S1��c�I��u,����������?>J:����2N�4zH�����9���ʕ+���~H�@I�������`ц�=&a�b7�G�����aO���\�Y;�����
P��3�o�=n����K�n�Eܮ�|����˩��s�ʙ x���O=eƌ�����J�
�F�$Q�N4�{8`�#�R}��8Э_�~h�2=��l�/�j:���iƃz��daEU�:+�jo�����af�w��ۻ�DX����l���F�ٽ�<v[�A<��:Z���hՐ�FzD�����C'�h�*\���1�c����sKg`�g�"��mJs�*���� ��%S@B.�4�JIE稚"$�J���G&Z�
������JD��2�U)d�0v��|�c�t\��|����;vlee%�D��ݻ9��S	K
���a�2K��)h*>�[��wT5��n3���g5��G>��J���B��������@��r�l����jhh@3������)S�us�-����~;��a�n�r�����s���1~�z`DD� �-�	[�_��=�����0��ը00@� +� �;��j������d�L�.�iV]]���c�1Xmi�ԩ�ƍ�&TUe}�	 ��y�Tɟ<���)�Tbe�t��a���T)��T�Y��r�1ǜzꩴb2�|����*g	 *��u��>��\&��"Tbp�h]��ic��n7���G��S�Y���ה�a��4��%)��N�e�^2*�;c�ze�bv"~�T/�Y�3=��@K)�'C�3��I�S�Ng�ڸ�ϑ�$4�Ųz�Ss�#��;w6�Qs�q;^wٴi�*W<Y����+N��R��6*4S�u���#,��H;��\�cP�V?�.0ƹ[�a.@>�_5:�7/�Qz*���;��������J���;[����T��ٌ�PS�r>��֬YǱ�Q*�A���[�}�]�a.�Ui��-\��nes���"d)h���\�G�[��ZZ[�����k������~�̙��L�:``�I�Q1t���vڐ:���%�\|�9gG"���x�d�W�s�p���,�ЋD��ׯ_�hѲe��~�m�̇$��y����A#�����C_"D�#t_�ziy�L*MG݅%�����y��Ka1lp��/��bӽ���1dZ�θ�s��y'��:b��)2PX���K&L<��؏��X4�M�V[�OU�ͅ��pQ[[������N';�@{t�;�������儘DN��;�)�X�>��]Y��OF>�L����䭪��� Q�ܽbA�gwi��� �Zb1lL��r�{Q�"$�h�+�<|���0=��b�� I�%0��PQqI��yn�7DH!�Eĵ:Ci��F�G�Ia2%%q#�qǜ�fE��Y�.��C��y�0DIi)0.���ū�[�A� �q��T����Y�f~�[���������1£V�3��0���'7gΜ����+���zԠD��uQ/]��	.�3��(���^Du|v��po�m�u`���.��{i"�s�{�p
#"�x��gO;�/��K�뮻�O>amG�PV��v)! Y�ӄ,X�������@W@��&w��u��H��dS� � -VƤ�������q����ʶ�,�B������A6o�L5y��qe G;�HA��b�A�]l�
��=�'�c���1l��S"����B%\�jkkG���N��'���(l�u������#%#���ѫ���i۶m��V��z@��>5���3g�֭:t�������b����J���ENZGT�m�4���\ y=e��)����ךJ�b���t*�����%g�{NIq��]���>��m�d���ˍ�I�K'�*	�����ّ�����F���mmm�t�D��Jg ��38���>7�իW766JBp��y������w��"rX�$X�s�J+qEOcC���H}|�_���d�榦V K�+S+�R�*�'B7/��3�<��O�%������x�_��(2��#8���k��+�Rr�XE~��6c���m����O?3f��ISƌ7q⤡C���WYY����ȅ��P����f�	�����H$�����iӦ�k׮[�q�z�ڵ˹�sDzƟ}(=���#��Np�l�����	&h�N1m���Xn������l:'��i2#	����-�X����٦<����MP�4T�-����<h�
����vGG&۠A�Dk ��}� Pc��h��SBv�u��<׾�#�A��Х���l����&$fUR���%�|�f�D�(��.-+f �!�N�/�Ø0��eSK����$��Q3%Bڦd����vG[g,��_T��i��C�HL��;E���vP�T2c*}s�X�<�	t��s��lI,H�*��r���p0&�ZX*�3�;�L�;v,]7���D<B�-�/�B'�P�BĻ_���[p`G����C�R�L�8��p�UVT`o�F:�Ta� 	`�;�ėZ.�σ���� 1��@V�|�S�?��\
ύOcz��S
B2�Pg�0��(Tne��!5�5@��^q�]wM�:�r��Ǐ���(z�˲?I�1��@�d���;w���G|X�1*^Rf�Y��'p�����R>b��xf
�A�
nz9�p&�,4T��2 �iH㽤Hys3��uf� �5����)���X4�c��.��F�E��2%5�в39�Qy�!(L����Ճ���ꢦ@�
Il���C���_�w�y�r+V� ��٬Ty���W���xG�9v�h��C*�u���ŧ�SlO>�@M6Vz`!���FnX�i��]R���I$�Ƴv*-����&����
dD�y��SHG�G�VTz� .%V�s����+~!�	����n�z��TD���o�|��3,JMi�a\���jʔ)�]w�[��ZZ��š3�p@N0�8�q�����;�+#��ga_9�5���)��7oާ�~j�D9�������n�S�[�5s!j~�8�����ٹ��;���y�駟���JT���DX�ef�qA�i>�裻�{���O?��k�͓�m��aQ:2�NÑ}�����S\C�2]�h�ٌ/'��_��]�d<�l�z�))	�4x ���&O������"�1d��X��z`�$~���s���۷/�di[[sS��;	����6�Tb�����'BG�#���ҡ_8��L����p+���8�U�)�r)Z�u�����l7�� �-��˘���L6$���I�d2��	����9�e�~���Js������(��и}���Р���X��EU���9�I�����^_`��Xx5�k�:�,9_���nWk	On�{�r���.$M��O�B���cN�DJ`���������F%gHɕ�GE%*g�?��e�}�na������\�>z%	�v��9�r&�����җ�T;h�
�	�"�~�����7|*�n���ǟp���DkU�7���Q(��60��`Ӄ�	����ꫯ��1����3�Rs	ׂ�KE�D�)Џ�d�yx���	Е�b����2�����8\T,_�F�Ej�����	5n�6
G���� T1Gy�.ÑbK���gt�N�E��Uo ��j'�>��[o�\����{��#PR��O$B��mڴ	� W=��c��~{}}=`7��Ix�ȊI:�����M?�oT�Ǘ$���4`k[8� �Dp,�@��--s�զ��pI`6Y��9���p/
��~��d��رK������
���&�:��5_�
U؇F�����K�|n�Pjjj�qALv#������---����x�݁����I��pʲ��q��O�?�>X�=��x���_��|��ŋ=�aÇH��J�+.=455�FX�'�x":J�Z�Z4����\e��Z����HG��#6�[�N�*����86�\V��|,��>a���3����ǆ#9�W�SI�)&���4i�,�kǎm��m��g�yjw�N�Z-^���d�ԩg�qz(X��	��pYq"�1�1��mێ?<?���()|�7��5�+�ª�� �X.{KK�#�<��+�tv�$з0r*�J̠S��z��G|�LmR4�h��z���yGe��3�"R�Gz[I�i|����?`���n�j՚+��`�|A�����p�(\��tqڪ(�s�������$m���,��x��J�~�z<�>O"t�_�=W�C��!��$"Rq!U	�+�ngU���-%�\
I
�KBh�pn|}~�T��RPOB�/8x�`�GWiQ��ǟx�=��޽]��2�+��l�9#-��t%�fo��L=tg�V�W�8�S�K������r��6dȠ\�]^Q�ud�c~$���8q"�~��	G��dJ�E��@�>�xl,�yx�*_���&�T�p��Z�k��f�t���x��(J�L:/p��HJKKkՁ*��Ԥ3i����!2�ר�L��xZ���o�tn����z�t�M�p��+j0ʥe�W_}�e_��J�.������e^)E��'$0IB�ܮD2�ˤ}~O:/.)�V�>��p�Q��.H&4���d2�G}��_���k�=z4S#�$�ⴝ��A|���Y���r����7�| O]V�5v�9��Ie��*̌6h�:yU���3�T� J.���Q����ʒΉ�W�X�(,l�T kա;���ꦇ,t�T�SB�R"�����"���_x���1��jr�ʋ/���� t�p�B ;:�Tu�}��;G���ikwZ��K�K��/��]a:�DO<�SD�r�1m�b��g���=б�Zl�/o�}Kˀ���Ç~��}�Ne�mۆ�P���N��9۷o���z������Ɵ�p�{�y���hxLR)��u�ց�_��xpi�"�h��ߪ"z��	I���ml�j�X�W�^�t)W-��[[�_���`�ߘ4��\w�7�;��7�xw�vG�Y^^�A�X���3g������b�������-� � ���y�a����+.�t͚5x�ݻw�����k�2{U�lN\��uҜfϞ�����ۊ�J�J�|M�����3�o�U�&��nȐ!ǌ��K#F���uu�TElq�|�K�Ϙ1���m�?�SO=�̇��>gZ���"~W��s)Oc�i��6����ߑ�B�5�������>Uc��0�ّ�ta+�'��d�pz��1�[Φ3>l�L���1��Y9Z.�%���X�Q�t@.�m��>�A�{M�6�=��Ɋ�[�JF��-lc��'T�A�ɨ�d�iP�{��K��DhR.?[�����3���3:��IG�O>����]�P��d�z�Z��b�dنr�(Af��w4��`P#� ���Q��W��6�Ie2���'�x�W^ѯy[[G0�I�r8��u�X,J���D{{�!�*fFE�I���tz�}$�!�R9*;�l�J0/�����Fxܡ����@z@���J��@�ׯ_��>,R��.r��`߀?$J�}Z�8�T�Q�E�Q�e��p�[�>����׍�gS�\EY�۔`�L������+Q��_*����S�R��Ĉ��e)W���a󷺌�!��"Z�4\�U�m�JJC�z*�*--.)-�� ],����PЏ���	Wlg�̮Y@�f����pM���{�~˘1c��j`";��X&* ������+J�j�����@��=�LCc�ǝϲ��ny�t����"]�J��,T>�|����$�҅^��'˹�u~|C�҈Ϗ5�)@L[g�KgT��	��&~�����;�Bɚ�tx!�Xj��i�ڵ��|@Lo�)��6����8�B��.)�-:��?̄!��u����v�3��!m����|j�9�x�b	�𓤅�/&���@����Ҙ<��b�O�l˅�"	UQ��ï2m��B��6�y/�ɞ-�0�N��$�`acy��G/��f7�0�RQgVQQ�ۚ ��2�X�w�}���V�O�]u��ԝ�_hc2��)Ҁf���s���S?{��w���;�Jb2�KU��0��)�3����D������N=�T
����c9���R`�H���R�ښ���T�%��[���拡qJ�^�����'�3j�2��%S�ʩd��k��3q�x=�H�=��QH6��.��ݬ��񠋒�U�5���_��*�{��ux=�t&���/�|�����c��p�ō]2o3��v�1d;-������ �����Ӈ�a�oGc��c.���HVMilN�\ZA��
�XE�G�AL�d�-�&�;Ovm ���n�l"�s�+�/�Qu��+!m�<Я��+��ʒo
"��jMO��}
(�<,}��J.�+������[���m�e��c�29ز�����������]�M�l�2T�NG�3����vͰQ*�F"֯[����mu��׿�'���8�O�U2l$�͞={�O��㱎����/b礘���x���m���D2�-IT�l��������}�{�2���I�T��>�r���&3!�=v�ۇ���F,C�켒m����7>�ϦǕ��O����W�D(?���!���ɀ�M˽n��W_}e���Au��xq�3<.կ_�Xc��i�/��!����piI)ڝJ'Lɤ��޽�������ږ[�~�d�@I�H�3�*`�7�x���+�r����ކ�O���G�q��M�×P-���¢��b�p��(��ά$��P��n��\�N��ɬ� ��2��?���-ۊ�K)L�:�ʨ!��H4��Qr�[:�!��3]����Ď,���-]/�W$0��`�z	�����xQ���B�K 7�3CC|n�$H�ylK?1�D��ȋ�H�F�2�v�,+�Xju8�Ӟ��ӧ�Sю�g�Ν��Nqq1(�8ەJտڛM:$����ؑs��&m�b�%� z���]:]�q����]�vQCs ���0x���� ܘ*��Q�>:�ԱO�Ck[3�ٖ��`A�H��S�W�Cm(�A��+���֭[�bȏ��(�fU�%M')bJh�X�!zw��V��x��d��:�lق�������4��G%�|%X�ؿl���y�늋Aذ�`�v�E%�%�0�W��V!WYo����i�� ��'����Je�RT����J��-E}���J��am����cb�`�Y�8���P9�`k�s����T�����b@�{8���H!�1���fV��J�r<�J�,uV$�pR�ܘ��͔0a8�ފ�dD:¹�.��bq��pBZ$�l޺�������f���z��\:�q����Ď� ����Y8�,��C�y�M�Ee�p��$��}VD����2�/��-8��m���4i��X�}��$X��N�e�f9�������.�W�q�b'p����Ϟ<�k_��R�3v��Qi!��6���z�l�Ǖo�{�y����[���3�^��Q0�YBN��CԥU��R۱s�������2eJ(\�����H$U���!�Ve���t*�q�ga���ز}g��NX.��%��4�Qܜ��;���X$��F���"����E'�0{�	�-�ʤ�^���� 4+\$QUL���{J���&=.�
hhn�R����'�n�l��d:e�.]\�2�
90��X���+��.���\�n��q��v$�9|�0|xɰa��Ɇ��2#F�ܾ}{sssmm��'�<e���755}���W^��]�0q�(��UV[k�w�.����J��UU�,�Y�+��H�tVg��5�܇�6;�������I����!N$+��z�O)g�T2�g:��
rO��z���b��X�^���F6�~��z4�֧њ*@ì��$?:�`�RK��+�����񁕍���)��x566����a����v�0�/ƆI�h�-�2 z?�Bح=i�m/��.�M����[ZZ�/_�E)X����ڊ{i�M��ۦ�E�GD%�.�����g+W�����G�A�n> f]�N�2Q��O���_��g�E��:����y�vv�j���º�L�b�%��/�K*���L%�*�s�l���o�v��;Čë����k1FC{��[(��m�f���0	?��ա:�E�+�-�㔗�O����Y����9���Q��콲�=6Ĺ=:�y<�|�G֬Y7f̘����"t�����à��z��SO9-饗�Ν���|�n=D�	g�a�Q]�Q5�g�yq٧�ĴF�V��9�KB���l��@{$F��.[���ޣ��N�^9@X{��e�b��n��[d��R-U:��lco̡��>)�D���e�G鋘��p�L�Y(D�E�t����=y���:۶a;�5��%�REx�.�n3�%��D�D��X"��L7"���x��X�i\8 �uޝ{u!Ix���BsmΝY�K39��$B<����3]��|V/�W�gr*��`����[oűw��*���L$�c�S�Ҏ��pqg�{�}�m�[�j���k90��E���8b[����q�~��7�|�^:x�`�������W,[	S[[{�'���4�������ګ�=�ȓ��q���g�f����R�dȷm���_xv�����m�,YZ;p��Ν�[��p�VW��߲E��uu8��K�Jkjj mc]�8z?�ty*)jX��"��&m��د�Q���D&`�i�����/����/. ��>RJ^��Dn�D�����^�ň�b�={��Ы Y��X�=#��,��E�ߔ�N�����$�Chzw�5�o����'N.�ׯ_")��@BwLoP�Or��&��*5ȭ�� ��M�*PDLBp�Z8L�gZ�"i�3R3^Yki�5g8u�GC�i����AGT�n�Y�2]I�b�Ad�3������]������ɠ}V̵���衇,XP^^�+�p"��8�D�AY�8D���;�	J�=��Q8��[S��U�,�0�|o�b�0O��l:�M�5��uqa]s���6�v'b�@�Pi=�I�FX݊]g}>��� B|^ъT����b**蔹>���4�@�޽{޼y���`�K��f��E2c�Fyy	s��(J��n��X���j-(��c\���y��k\�\k�%K���r>���$��V8?c3$N$����m��DGO'�Q�|��u��Gծ��:5Q������S�[�,�����Nn�cU�V��~�e8w�^Y���D�>��:~��<ի��uK0�Y��5k���عk�7\��%t(�""g������x���~�����%�s>��,���z&k���#ͬ�M�5y�w��L�f�};ԏXA;;::@<�L�2l؈XL��46�X��={ZL�'��z�I�OGQR��|:,N�7ޘ�ɤf�p���,\���f`]����-�l���
�ojhDˇ��~��-h�5�m�"�gUy��2�E��uZE�4�8ّ
d
�%�(�M��<^3�Ȧ��렐��@������uk7�/^YUZ]=�mv45� E�fs�}V5��Epq{l\JI�춣9����7w5�L�[�~��#��AN:i6~�������e��=`׸��;X�SI���7vuua��ƻ%9�{.^���b�yF�L��)ݮ����@�H<hp��tc��z��X����u:�8�	1EA�(w���V�ݷLd/扎v`��6�����{�O�/J�B/3�ˋ��)g��s+sN3t)� p/���Ag3��j��p9kϺ���2H?��Ӆ��	��O�R&�����֙��z��%��#��]�g�� kJ�w�"��ߒ��-,#�+�Fk{˖z����B���D�SUB�)9D��W��GȎ��i��3N�aX���!]p���=���<�G;�#Y��w0o~��م��p{c�-�3i�	�=�G���;5�tj+�K���ϙ9�N�jf�_��ڽ^��r��>�-�[�n���;�o��3gNyy)�����:��������?�O��k٦���)�!2��	=�?�g���� d�6K��u�"h�ڼ}�N���z}�"J�1���e�>�� R���`5'AQ��?^�Q�֍�x$��U��o�I$��
� k׮e۶���;v�TB!m$>U�#���PA/Z����ufɊ���Ao�:�C@��/��Y�B:[�W]�԰�Y=�[Q>íA[�f����ς��[3��3R�uQ�����|����퍍".����WIQqyy9>�ÀLl��d*.�υz�{�iz{�:�1t"�����u�����������:��N����5����� �fLh+&9�����S�� ��C߬�Y�He��op�<d���
��~�K����es�.
EН�G�!��uIPi�as=N���/�w)b��T:g ]��Y\H���dPI�.�G'��I���ȑ��G�c��N�LB�뜇�ֺ�ܲ�!��[P!�ö{�������*[O�ǜ�[��]`v��ҠfV7��{%���>����G_��{���Q���W��y����	�CH�����h!7{:���$��i�M%��ӈF,&}���cz�"��~���>��UUU--M���2Θ��	�Sv0�7\~0������Y�s$7#���I��J�-�a�\�I�j$*����I/��^c@M?\��I���E�^*�jf.zmv>�W�����+YI9�� �%E�ϝN�$`��$�=��D�;�,ԩ4��B���L��"�^�ޓ�S<&��r���5Ȧ��p�=Fj��S<0�4Ad>&��R��D"1�?�Ԝ���8��H��"��;T�!p���v������1&��K0�Rɂ��C4�l�Ӭ}�����X9u����0�k��"���3�� �)��c>�XVV&��J���݃��u��Bĵ,uJ�!]%T�a��B�+�M"k��Y���up�:�p�)�-��Ǆv�id�;���֪�$��E�r�I͂���(ANԃ��:�<XD{�^�T�
Jh��vZL��u�������a��p�2��{���lF�Z�vsu{.��{o�ۣ�l�`�w��q�����E:ng�yE��3�(p?�:��g���?�qiC�e��=`� ��im�Ƹ�ւ6��p�����n����o�`�RW f^"���A)-����rϞ�fC�*|^��0��J.J�_^��eD����Ȳ4+���o/��}�^f�zf�̀��a`a�!lcl#�e�B^cDX�� �
	12�����g�^���kͪ���3�������?�|�eVVvuu�t���|y�]����;���� �9�U��]���c������\>�l*���((��riii)�ӆ=�5��K�S�˖i��
S��/��d&il���1ܫ���v8�����E�� d(���ATT�&�Y��X��}�� �.�u�\��Jx|�R��r�YEL^��\=/ssZ�x͔Ǎۃ�҂�^L���������C�WF"�h��n�n%_���4��e�kM2�(%�w=bSO�*��Z;�����̖�4��Gz�U��ނ
����:�;W�@�k���h;� �#��P�d.�����~�=�d�&m�Z܉'��Az���ȱ�������T�#kd��u)3��}�O.c_���7\\;������ì�o]���R��@馴�~�#AB��һ�Vl65��.�.2)3\��Ƙ1��v��|��!Jk�2�R^ ��5/�R(���?���c���!4VY֤��z��%��힙��ZX���;w�H �]z��A�X9z��cGN�:u��1A��e�'9�O�7�������/���Y���v���u=��W穤L�	��W��x��.٣�M1�O��):�r�����j�irRꖡi��잞�S�E���=ll6p0$�|�\(I��ȉ���r��8� ���i$�G��5C�E� j��j�Y��ժs���9`ܫ.s5V�DI!�)I�R�s*���\��q/B�!l+�����c�f�Az@�{�,���RF���r}8:�C#��M�q�8��P��������&|�5�r��D�]���xg��y�g�t��Ȁ�Ȭ?�u�ځ��V*5��ݰnJkU5�ٵ/+�˭��2�OyǙN|��}gx)i���8r������K����J�������0��m@�� �t:bU�P���9���;oG
�
�r�n��+�5�t�h:����Q�K:��^I�/ʉ��2��؏��<�\X��\�C��y�w�1�ܭR���-�bMI����}���%��|��ǎ3qo;adE�����?R4�\�����4�z<�%Y�x_��� ġ���^��ȑ#�o�7���'����P��I��	�X����k����������V,�H#��h���b[,�{I��a�lIKe�e-Ŗ��������<�3$>���z~�f��v�o7[.F/��S�����TӤ�bF)�i���!�.h�0
E͎�؞)�!	CK�b���Xd��a�i���a��X��@T9S�w8,���@Z�D	k;�zna&xr��΃�۱A���-$����XrcDND|��	���%�(�Nwv)�X;����z��] ���
9�j�c7�m��b"z��p�$��fS9�U"��W�w�𕹘��Ƙl`ee���8�A��`&�x*|�����#`#�E�.j`��3K �
���`��!����>��T*�7�_[V�~]��q��EC�/��T��qJ��R�I\�A<5�,��'<-W[�r
��"OW$���p��v{`�r;�/�^�;c���t����\�j�?����eg	�B�f��QbZA��oF`D9S���W��	�����c��'���
<�t+h[�I��phߪ��BA�����(�9(��"�ݬ�ږ%��*A��QU;�?�>�;!N|�[���-�*WCtq��Q,���Q!w5T�D�a���*}E����������������z��sQ��4l	j#C,A�F�E; i5�D��fd)�vU�;��nGb8����8����H��SP]���FF� a(-q⑀PU�&y+]`�݂�H]��mDk�밖
���p�`�),EJS��!�-l��(AQ�̙yA�I�)S�Nw]X��K����At���D	�L$�q�����F�A2�i�x��Pf9#&
#�����PK`���i{PNë\PC�dqEAW
��"B��
^��'���v�)Gޤw_�C��¢��"zE�*A�n����1�,��w���id9���I"�ll��9[�c&j$s�6�i�yc[��g���Ƌ���.�J����t�7�	u��X?����.���� F� �;]�3_�O�j��{��k���_N�y�}{||��l� �����UI~��#� u�cś�'۾�zey1�������/��X�H�KW�7Ɔ�dtW�����Q���3���G	�l@9#Z�e4d�?�P>��C1O�Y��hxA�d��;A������ޙ,���#]g��8����g�'����	�0�1���jHYjf�-����s1r�Aŋ����)Qc�i�,Ô%�2���Z��*q��&�:~�r0�mT��fTPQ��0�D�?C�=�>�n����	���}�����.r�x0�ccc�i�牉),���9 ������� ������G���ۿ�߭�nT��k�&����M���nK�0�&kI&"U��|�۷^z�7$w�P�aSEcK2���h�f��h�˺&��_$��v��u��I���!5��m&z��;E�~��y���W9�qUS�H/��5{���$�{ݏ�\�g�S��ӡ���G*��N�k� ܇l�mS�̸�%�'1[��jM�c�^dq����:�O��	�J��3{�R���8G'J�='���[�P���P*����`ve��0�vC!���FR31Z}�1
9L6��~\��/.�U�2�.���<[5V����쯁�����dyK9̎�Զ\z�/��)�)	ށ͂�� �Q�V�.)d5�R? ����q��Ȅ7�#�I@/�JĞY��Ը=�����T�^�ъ�T�����{<�{��K�};7,�r}���@h)�?�ccU��&����ěI��n����/��/~��ϺN�P�}����݅�����ƪ�#�'�֠�N5B��K͎S���n*�O��P&�����L�w�3�p&лG9J��,XDC���5��L�}.�x��#L`gc��v���֛NRx�ܙ�JpN���7��q�|>?11!�<�oq_Pa@B�uџS%����ᑟ���p��|��IpOP��M�(� �}@�?b����&�E\��8}q���	��=�!n� CCs�+����i���� ]zj�J�ON��.5ř[|rwQ�[��3{`�_��$�Geubi!uB%z�������m�㻦�!H^��RS���W�jC�|_７�
�^{��?����he1�,ϸ�R-��T�3"�3��!�=�o ���g��J���5>�&�[e�L03�'��\��C��e��E���&B�TJ�,c6�'���"WadP�hb;��R��Z���V=\�����ƷFN�C~���ÚV�� �uK�{��d�X��r�֭�ׯ�����O?-�������Q��������!$>�=���'��c��\�4Y�����26�x0=n�޴�7�N#n5����4�Y*���i@Mr�߀��A��7ư��OZ��r��ƽRAqŧeF9{�����^����=^v��[���V���T��r��w�S�(��8�WŌ4>�J��iώ[�M��Կ����Ą� ,��+��N��,4\����h��:JRyq{ L"������_1��\��f>�$>����"�(S���|j�}�_�ϰ�1�Z3�6G�
�	o,T �S�9�4\��XJG����C��6D��? �ǻI	�ҕ�Xe�4���i��5*į)��cI��	̧O�>|�p�V��=� ��`�,j�ՇL�R�n��u�zVf�l:J�+�;I�K�O���x�7n0���ܪ�jh��;��M*��{Q�T�w�$��?|?��C�r��kD���˹�vk�P(�����g���������G>T.W-[����_��o��o��������a�E�X�����$�-۔�<@����k��z۴�2�x�Û68���(30��*3�E@ �D��Z�T�"�n��j�UJ���,�l8�YLB��Qs�T�>��'���D0U�����C����s@@�f���>���]��-:l��gffo�����`�������p�(����t'��X����r����	�(s���v�}�U=����������#v���NYܨG6��
(� <@ÿp����I�*���T��#9j�W�7ؖ�G��ZRm��o�i��)I�%�7W�h[I����}�R��l»�;!�.�w��?�S��k�(�R����4�C�NLL@�@}�S�����'O3��p~F�㲢���TU���S&�P�O�&�>S�
w�Vd!!�#P+A\V��z�������ݵ�5�);e��ً\���9�m;�0�|���@�������E�=bz��|��Ѡ*b��(#�_��41�s�;xp��ۘ���_��ח��?�Qn�
�쬄^f���aͰ?��j�jim�����Ye!&o�b����b�����HT��3seF˔�'�~�	�z`�n���d׵1h� 	��L��-����B�4L�A;��5&�%F)��$q��.���v�B�Zr�^���{b�a�";9I�t��$�g�%'�|��ӧO��o~�*f�X�þ�==�f�ڶ�
r?��Ap���X[]��2�ZZ�;� sZ����N��_��u��C
#������
`�EmPZ2zd�����j�C�:��I�#1���g��<훶�UD1*	��,ʄ��[�ʽyd�=rq���G���j���Z��A��k�=��� xWV�._�,aۖ�EYv�l�;�N�|���5����O��~4ն��VJ��x�]������(#��j��#�k�9�h�B9tQ}}�Z-�y����,s�?<!��S}�.�ݛ=�Ǝ�a�lI2�����9��&�hG�,�`���a�D3�ڎMIt�^~��K/��>��ll��+��?������3�����+�B�=�8{�C���DE��o��m#j���mB"JF ����	�a��։�ZO���d޴��.󕋹9Z�-�H�nvdc0bT�Q��{�r�׭�יM+NC-�?0��k$F ��0�f$��	b&�E�.�X�=�3}q���e�0�\�B�����T5��=W	Q�^�k���Zxuɾ�*���P#E*��D���~�/n�V��pw�n����D���^���p
��	�~��1�:�Аi��p2�+D���b��q-[t��ژ<4:m�4|�uۧ�v�鵔���`�:~���x�a���F��^�4<Q+������=v�Ȯ�<��G8p�=��]�y�����Xٞ����q��δo���U:���m2==��?���?�<�����W���_��_�?��:1(Pɏ�;'��Ϟ=������ca�K`)�����n�!N�#p@C� P��{�0E>�n$��YH�V�Pˋ��Vl˘��y'Z���� L��/W|p Jm|��m�J~��f>������X �=yV�,!:��a9�	ps�X(��-|X*�������I���f!��X{��sT��2��F���e�����
�):�Dd{ItIR�O|��N �p�С��D�w��RME���=�Q�����H@14��T�'��ggJ5A��v�Fq��Ɩ�<f��6"M�X�U�`N3���
�6N$I�9`�9���?|���qd2L������W6��;�ծ���`�����8{
�����X�*������R�`9H���e�n�·���T*�y}m��!Sp�T��m�,pH������|�	^ 	�=L�S�N����sL�$oT���+�zh�⻳��"�6��b��ÈBMr��p��@��ρJٺ�>��2�\2���|�&�H8w�^���u���w��yi���ۍ�����K������ E����&���Z�D��Ǚ����o�y���s�?�����}���:P�pú&kLoe��!�=�!�Y��Ԛ�_$5�`"U���(!���<�;[[_���Z�v��1�a/!g�E��2m2ވi����]:���T&?6g���@H�|�]�ޅ�Xje���C8�3?zJ��e�M���l5���?�����کǏ�V�����?�����������KD!��%����W[�jJk���m6=�t���.Y����������Ic-ԍ��� "b��.��)������ƌ�D�;̞�$�NՉN���H>��$t��	_}��3�<�裧�]�������ə�$�Nb^wq�s�f�- q�!m��'Z:!L:ݱ-G�OL�)�B�ks���#��]ZZ����ޤ������$�[�d��<��Ga�3�%h�&Qd�sL�o_�|k��#G6���n/�C�DDS2���l�||�Ղ����\��w�EێR�ck�e���!֌� �Ҵ�c9E;��!XҔ�=�m
*z�V������
�� �g�z�d�h�*
�0P��� `x��.8ݤDì�h���f���+`�F��S���MѼ����v�D�Beu��X���4҉�q`��_�6�fbb�:����^I(E*'jg-�c�;�|B̒���"*]�_��z1G�������GtӸu�7���R[�j�2Y���
�������,���R��,W+���cu�+xyMf��g�{+��Ï�jkVQ�B���K)U���k@i��9鬺2Be��9x����q�"�ټ�j'=^*ü&{�b���,��_Iv	Z��N�c��a��S�_��/��_�/t�a��J�2�����+oT����O�8���8���	v�Zq��Ճ�������s�9���x��L'Q����R�M]�d��c����@R� ��K�0;Sǲ��5�E��XX__ǿO=�Tul왳Ou�]~��F��lR����l�����n����_��Y����Ng�TF��C�h#����C=�K����|�1�:�`����{�R���į�����O=��vmK�������������1a�O_�ܳ�c8�j��y�@�;�#R�BQ��h�}�M�&4�c!^��,Y�)MyF�,Z��� ����,yR+d;3N�ʴ2�7�$g�h�(%�{�h7[o����ډ����͗��#=	$�;&D`�yƟCø9�5V�͖��26�q�PP"R���<��^���%+0��
�d�5	rhu��,�J4�J��N�e1��#ҥ4';酂8�%s��
j�E�����ky�ǀ��g�hY�X�;��H4 ��H�XO��24�q(ؤMM߱xc�I���QSFo��N���DSѣG�rP������%�ˉF�$v[ͦc#;N,��0M���W+�@�)߉�"P��1Ɗ"@Oy+蔊�Z��~��i;��|�����}��Q�Kn�X(:8A��)Kp
�t{�*2��k������@͠W�5�m�N��U8��t��*K�ڵk�C333����[\���f���T���BbH3==��+��ze?VM���cccǏ��������i!:�s�����y���R����!5N�g����cR�0s�2����vd���w�;�m�AY���a^Hl�Д~z��l�"SF%-��Y��n�#�|d?��%�`���c��RU2���_�˯}���Esu�ת?�}x���MNN�
yh7��#��.Gu4�SM��=���2�5�̍ק�D�d�� KP���C�&�S{[�mn�Q~�lR�mf�?}�4U�6����1*�6L�Pa7n���W����z���xk9� �H�ֶ�UPm���V��v{�.�T*�hr�;�	�k��f���#��_��}��4	�����g��?����ܥ7�]�75�SUO���p�n/�e�L}�Ɵ���W�¾�u��D��ȼ��w@�_4ݦ}�هM���a�'�
��������+r@��}�L]46���9?�����0�L�cG9r_�s�j�bK���Ss�4KLӲz�X\�e���S-٬F�g�z���i7����D7U2��DN��tKvV���R�P��i?\c��u'���)?�#�d�N�݉������R�vtj�L8�!�#3.�W�����[�n�Sp������%�ϔ����tP����6]|%Nqe�uʥ*Ss�A�MX������Ǉ�o�^\�s�K����;��` ��51�Ϲ�]�$��&��i���L��p����7�i��è���_����ٳ�n�V�ܽ{�����/}�;~�S�-#G�p���gL,Х��Ϙ�Ű�^�V+q�\.s����1����y$�I��Tz�srX`����z��E��\)����p�C��X���d:6�T�i61?���2��{��v��g<�BhP�kƿ�NіXK��`��jB ?-n�ޜ��s{0d� /����B�SOw�dv�X��_L���o�U'1����j��5R� �J%�R�ЀKB6�{����:W�Z�)]H���-� ]�luz���/|�j�?w������j��]�0�~φ�g�Ը���*��*[���������6H����j&�)�L�]��$��B�_����6m+
B�Tt;��-&�aRD���nX�u<�O�A��l�
�R����畕Jy�Z4)�4��R��[f�H愿�@h�������}�c�b�ۏp�=ll�1��V�=y��cG��B#�7Ͻ������y�k�j���HD6�J&"Q-�w�-�d�N�Od��;��AH�z�|0F{X��c�/S��7�u�zЋ+%J���-|c����8H"X������E��&7��yI,x�(��\���р-xwa?OLL�t���`#P�&{3K-(|�Y�Z>
�����U��qe�G@(\&�w���k[�RŴH�bfq/��&���M�"I4�%�Ad;F���ego�N�d˶RJ��v����Ї>|��6�MS��z� �r��:���5��V&�0<��z^�ܼ>�Vo����N��L�L9}擟����4�.�L�<66���Ǟ|��0v/�->�����O?w�ʕ�����bc}�Knޜ���p�����G־3P��?��@��*:*XL2s�ԩ_��_>}����p��'���������E��QZ/��o�!U�h��&�adi�'N�����q�	0�/.�;�2�u����o��	+�
������׿��s��QV'mL�PB-]�v��G��� �I��.T��O"�)������=����!�����ׯ�Μ9����yI����5bTm��[�e���m"���p�٠��Ż�Ǐ!��W�y�Tu����¡��T%�)�%j���V��q����B�G���퀮Zx��������B�����Յ� ������X�wn�]o�Z�|	T��.U*��%�1	��U7lU�19C���$D�(���龔2T����L��o��֗��b�$N�Ȕ�f�z���#��U�Q��J�V�����3Dc: �N�rm.]�t��U�6�Ou򣐆�x�u)^f��B�ze�������ȏ`} ���[F:^��V������o���~��W5�n�z��fh��w�$7t�V'�7���iQ�^B�>�O��OK���H
D�'rlϊ�ִ�Q�Y"5�w���̚w'*j�0L��� �ž��Y���Q&R�Z�t�Fl6i��v6���Z��9F��$�̗�^�J��8Y�C�y���3�x�۷o_�����2�E�]�{عv��QS�8ba��vc���?v����
��
��(L\�.r"�ͨ+���#�R���iKr���nwwh���֙��pMO���O�$n���A<55���,�$�Xu|ui�ڕ��^~���<��������sżs����ǟ�Ƌ�"�7+����{n[��g���g>s��!����E� kU#^�L+E�K�Gy��ܸ;�Z-��,���_{e}}��_���p��Z�6.8��~�>���AJ���"��~zz�E!Ɛ�NI�S?�x�9,Ե����_��?�Ûs�(Pk�Shi�pr�H`�O<�ħ?�i<�P �L����y.�����vr�z�2��^{8����\�y\�z��<���`��:q���〩���`rߩ{S�-H�WU]L��t�p<-g�I�K:��=2l�o�(��했1n�@�������/��3Vu�LU��,lX����k���Z���U�����ꦦ�&��2D̎-�ST��}�W��I�Ž\�9%�SIz^}O������M��tiY�@��+�\!����vO0���9�4�յ���m��6vl���vd&/{�V�5V�q �7� c�,�|�KIw'��m� d ҡј4�����`�y�S���E�E��)~5�7+5��,A,�2 ȗ'�t�����xQ����V�R;�og����Ը}�����/��'�'��g�¤&Ap���k��v^t�I����7�|�+�G������K<����'�(q$p�d7ma��8x���<z�h�Ra��-C���j��Wө(=r{�R�2��a���t����F״�n;��E��N�vb���01�lڥ��ɓ�����4��6��\�+���M�N�����v�	Ú6�A�O2;9a���WϽ�Z�� ����4dO?�a\�}�5''�>��O<��s�,Kl�\�V�	���K��܍ۍȂ���ۖ���,����o�X���_GQ���m�ꢭ[,�~�~�g�����5
�3/�������kkk����*0�zcF|��w=�ܹs_��7�͎b����E�~H�T����"�Q��~���R��X�Ѝ�j����=���n�9tp���~{#�Z㵒h���c����;<�q>��M�T5�$UE�63�$�� �)v�mS$�A�E�~�b��a�T=��a
���&�T��#����3g� (��ƪl�ǂC���i@%`�)����|�T(����(�;ݶ�ka��3�I2l�`���ulF�����7���/c?���X$/���������ON�S�ݥe��ѣG.���_}��#��d�M�?66�tZ.��K'�1y�f�ڵkx�.���I2ǚk`d���SQ�D8�匹��N����bKһ��b�V*���j���.~��_��J� Q�,~x�]B��n�K��m-��?���m��������-�U��Y>�/q��I?��P�،��=z�/���V?f�v<cK��W��1?�R�g���x��6����`>�:mj�a��.��0�,'�Yd��h���PPY�(�	���X�h,--@U�b�g�C�ż��#��+3�PK~�!�2k��$9K5mS�bkQd��b$���E���e�0�Y�.���~�GV����w�<����ag����e���?�����a������SO=EFLD)7�<�`8K��������V}e�!����HD�}����Z���Ѭ%�T?j�T �����x?S�߯�l�r�K�b��m��n.�b�&Q<1YH{����~�+_�f�u]��VL
@��7��
q�	s'Gi�R�A���|������n{Y4��1�����i�7�� �j����������+׮�a�#�;��������u�(4��?��mvr`�z9G������>��<��3��Q�G�7^|�+q���[_�b�� >t�!8I�D�Ri`��a�d��?�`!�nia�6�+v�mH	H�����W���5��4[�ScO?�> ��^��l�����M7�����i�\9u��D�j����TR/z���-۴l�r>�s�g�ޅ��˹֝��~�ch&��Y�n�ip/ǹ�?`�u4ƙ�@"Y�䵇w��y��\���-�^~��7.�:��j����1D��@�Fe����@�X��X�|2���9ϫ�+����V �� E�֚夀;�T���,��A	��=å��7o�=|dvz��͛�q�=z�A���ݎ�:�[�����7������?DX	�%ŸNOO���)93�X4qB�Ѹx��O<q��A���W/�qJNR�NSw.�vH�W��&5�Yss�n�No6�F��<���[5%e�;�H{�C�c's���qqn+����~����ǻ�V�<#A[H���~n^r��d�[v���R}���׽�P�{vs�F�܍M�gg�Y��E�Ǧʕ1��ذ-�yN1_�a�+�&&��1rR����4���hֹ��,6����Z�gM�7�>�,eC�Q}e��۷nݺt����1��]�2O�tl���|&�B�b�+o%MMgH��|��
�T���t98{�}��G�L�2^)�t�����/�4�x��1P>�!��> r�R��o���E��'!W�p'�~a-޺u��v�U0m��"FQC#H��@O5m/�ex}��%fz��juzz�ȑ#�3�_�	��s�ıɩ������j���F�^grr||z���7�(�sy?HT5�����	x���Zr�����ك�f %��ݼ�Ƿ��n�%ú�� ~�![��:������ݹ{��Xck;"�Kd��������pWlN.az��kNMM=z��_q�NrD#Gv�B�g��6o���m�N����IRC�߄�(�2��n����͉����]i�8qdfz�(Z�A��Qa�W	j�,�vڰ�r0��7`�.c���R�j��X�6��A"^�ر�>�ccU�o�r�j��u����F���G}�ѫo\|��4躎U�H����2���e!*s�3P����`�"��q��M��T*~��=|p�_���⁄$��D7���$��֯Hai	�euXr� F�V���(�(�qL+#�j9_������������k:S&��1X>�f���'N�={��� `ҥK�y䑧Ξm6ج�,Ǐ��cO>�-s���W_�X��Y
G1-Q<-.�QZ][����ǲ�@����K/�������C	u�� Q����6�ȕРP�L�h
?HJk��i�dnm+G�dÊD���E��_1n{��%k�x��,����r���{k��m�m����q[��^s�P��2aQ��\niiI�bl穕�{�s����}Fҗ���}����W{o�I1!	�obb�>�R��h�ap�@�7��n����Ӳ������a\hj/GM7L�R��Ji7�G�$1��e�ǂؙ.�<��Ѱ$��
��|�r���	S
"���u���д���Uv�3e(Nf�Jv�c�%����@�σ�!�(Q�jYq$H�j�>��߽{{��A'[��h�{q�V�e�6�/mk�F���{�@�uؾ�W�S� 7�Yl4Z�O9a��m5a��物�fKҐ��MA�'~�=ѵ> ���B��	�2MiB"R\:�J���K���y�CG��|�+(�^y�����G��vu�j��Z�����#���n�Y���X6[�u���őF�)z�&�yF�c����kێ�lt��h'�����k�)۳����b�W��w��~���o^x9�9˱\/5�z�\g������"b2	�Nj"���4�Hʕ����Q��L(r�(iL�q�1%�6Z=����2pY����ۭ�N�91�,�)�IЈ����	�6^�I�dI��r���\�^ߠ�D�p�Z�TM���v"-�u�k+��������իo\�8;u�ٳO�ܺymea/��-|���3W�#۴B�<A��c�ӄ�E3f]�p0���*����B�W������GO��yn���n�����������DȮ�{'?>>Aْ�F��3�E�a��F*��-�2�2X$��5^{��ǿ��/E��^�[&E�M��:'lu�x,��+���86�G�MA<-[�:>셑mQ#�__�(y����|ќ��&�f�dL�6 ��X���&�k�A�z���+�K���<p`����,..���x�}��@�]���k.�
�|�gΜ9w��׾�5l�S�N]�z}umezz����ҹ*�(+�N�PJ�X�^�8C��<y�8�3 �]�a[Y̭�V �S9ߏ�*���>��R�pjG���1�@���X���6�ۣm��6�$�+.KM-�֘�O�\��p��0�����h�;�|�f����/;��k��ⶍ��б{�&B-qQ�v;��)�:���{�&���Mٺ��6���q&������Ւ8��wK�#��K:�y��תC��Զv���#�E1h�N�_��A3�$}��I�Bˏ�l�N�_[#���k�0z�N�٬�Q���ިw���+���_�A�X�^|���|�K���&=}�[�i��B�˝=��g�>�Zy�I���M+�����|҃�ilQ�U�8^��`�
0,��W_����yc�͡�G�%���l�E����QD�5����n�t��+���=�25A%%�Ydn��u>�/����^���Q���V������~�W/޸1�����[�M#&��H���d0+8���&t4�Y�����.YIlHe��w1Ò6Ę�����3:��~X�dz�=O!_�tz�	���Cj�����͛7O�<q��3�s�o޼�����s�2uQ��u���ߚ�6w�J}e��7�V]G�\l���	:�4�##�ó�K�#���jU�
؊��Nw��r��{�c�O���H�F7d�����`׵�L���� | (�t���������ql$}�ZVjX�#A{mバI`�zN��RZ��ه��8�	�ڪ��Z˼�}��e!f�嬸������Rm���6�>��ԛIEۭ�j�$���櫵������ߨb��A� p����5��Rwb

���7j�U�����\�r���'>���o]�ԛ�N�`�x/S7�{�H������Jc�̶ .I& LF[zDF2uC�X�N�Lu���ϩ	Nb	���$
i�bB��PN�@����7t�� �[��NK��Y<��� ?�Z'�w2z� l��� ���_"Q<g{���R�ф�t��a�������~�'~�'�����g���o;�>�`St���e�s�0\�R����Έ��ƍ�^�)q)\��!�0��j\s��I��ћD9v枾��V��H&C�|5��K���rt�s)a�b�8�_���J��#�]���+��A����$q�H ,M.*�;q����2g���7>�mbQ��������>�;ΩD��������a����\��}�p��O����oZ�7�o�Q���|c`��4����a�x;��1�� hPbI������a�Ԡ�5���W���������a�Aܺu+�⛹����b1��nVJt�ƵN���34}�/:+8N���lvs�1����j����ӧ�|�����?�ӕ��Ju��X�,.܁��=�p>'��}Z��xz�~�	c�l4Zݮ����M�T�.hrm�V�#�α{�Ab�y�LK���굫_����oܙ��4M�_g[�o�0�qA3�~YlB}��X��E��X��a?4	?����	�'���alc(�6�Y,B�;Ƚt�ۯ���Ea�<p�̙�gf&\�.�y��ka۴������N�<���x�v�T^YZ�{�f��1Q+����F�/�vb�X���<��F���,�1��jm��#�;.Q�ς�5�1rz�àKQ���/�ĩS�ʕ����q�ـ��#�i��&α-j�*`?.�M
�0�����)�UO%�c�7O��i��<V>�%!���ƪ�����=�/�,)�|�&��F�b�b�x
��Q&�8�R�שyS�:0s`�P����/]Xo���.��a,=�,Q�����6�(p_S�����ؤ;���33������ɉ�g�~juy��1�����Ņ;kˆ�S�qHwާ���".@n����	��,á޵�ֈ8:�(�ж<�+����[���R6�I���n�K�H�o�D���#@���+G	a!ʾ+���5 ��h��G|܄J������
�>�)�q����A����S���K\�!4���hU]�z���S'N�R�'X�?��?uŶ;N~��+�'C�6�DFࡥ2V�]������YXX`��O�"�����<l�.��u(�|��0q�<���}iw�����eN�
<�y}F�|)<p�Ze��$d��C͎w�i��ݐn������9뻁.��io�@j��m�)[�bɜ�]���l�V�L�d��C������(5l4�r��b�-�kN�жf��Ӥ��ɥ�&��Ց��w���*%�zg��۞SF�AS�{�,��*jAu�֡_Z�NL��t~�G�i��G��+׮J���������D~j|"?������������,�¾�N#k�)�m۰��B@dB�p����_���� �LBb��;����*�����c�Q�!K40��X��V}���~A���9��B����m�q��Db���W�<{W޼�q8x`��i�H�����y��B�c9�'�lp�B{��y9{~��{��oϣ�0�I��5��.��@��ڥ@��s��Jwu_�3��ֱ�m�;y��Ç�ZvbZ������U
�.O֪�N�
�V��{9��k�'Qz���J!�-�-��|M]v_Mc�j$8�K�y��~�_��ff��D����!-pʉ�ݩ������V�r�D34�B0��zl���8�B�a��+b�tڱ ��Z���v��&L�m��0��<��;�<��ѣǞ<���\�������ֵ:�#�]�"���ˈI���ݢ���]�.�Q�i4�������*�ۅK�n^9r`ƈ"=	�0���F�Cn�Q��.���}�����J5�:�0���k�v;��յ�����+�enbwHf%D�lxQ'zd}x�PD�0���f�k�zL�D)�Lw
y��6@gT�1���y�X�3��Re��`��i��N&D��H��"��&0'����m+�Ӣ�O���%�E,!z #]�%pX�ף*#Xێ�kw["9�@����LNB�$�c�OLqQ�W��e���y�Z�:/�Ç��N�T'N���$Y������6k���"6�����s�x��Ǐ���E�D�G)�"1)k6�ՠTe���M=N��X
B@��y�'p��pL@�ە�H���'a��2��K�l{�v��*���~��m<�lX�Z�ۙ���,1�i��u+����{ H�n{ ?�	e���_V�͛Wa�8x(n$�x�zV�X#�J��-�ދ�%�s�����k�pT�9���$ա��!K�+˓d���㳝Eeg�;!;��ob��㷚Iʈ���5g�A�sH�W�öZ�e(?�p�X�661�E�ؠ�Q�2͉�x�6�S]p�jja䯭/�&�cX1&;�C��CW���^';�Qfk���?�W'&&���61a��dq�UڟE/�ş���I/뭦���欭dC �w%����1�"��9׶R�n�����3'fg� 	�C��V�7�^C(P*�uD�4j����n0?�ҥKss�a�����{W �},4Ҁ�_9���&.��bز^D�O��Qs@&�T�f􄑖5Cp-{vz��� ��i��gzb�V(U�� l녯ݸ~=���B��)/NJ�Dd:Q{ԬG��v���0����#�GJ�J�162����F��#9r��ؙ�ko�e�uQ[��l&��Y�r�y�Fi&q q}���Q{���Z�n��Fji���(Nil����i�#��{��Z<0�z����)Ȩq����F��s�b�d�����(o���U�g���c�g�4�֝���6)�E��^tpR=�Z��Q*P�KyqUa��5*�q��j�7�k�a�;7��~MDr4K�h�!,���&U��)$��&h� �E�����)��S [ �-�2���ZI���{����b4�����c\|J��*�"5������}�F�^)���%A��7�c�y�vM�Ce]"�ǰ�
����~A���bzj�X��.��Rm���8�W]<��"�w�����u	*�����c�r�C1����6D��\�ƍ'O�|��ǹa+U��j@�[SSSKKKÈE2˩ѡ�|6� ���#$XizJ.5�a;�T-��W�jx�P�A�K*pُ�iw�D8.��+p8hg=2���Y��|FE\�ݠ����{��x ��/*	�U,S%"f��?0*���0\�d�k��\2�Vyp5*�ְ��p��rJ�)��R��8r���aJ~ȑ��5�P}fL�=_ۥƥq&�Ǩ)���s���w,�G7��,� *O��Ҧ'�?�я�:u"_,t;���rӊ�99 �|����+W�WV�����''(i��s��e�XϞKu��n�)� ���2A�W�L
�F=]��v����_x��W�]\qiEe���/��\;�tGiI>O�HR��F����Byt�����M�I��$�@��δ-��Ra��iZj�16w�&�y���s�>�8E�.����N�~����El�#G�OOO�JqM}}���/z�K�͛I��n�TW ��x��	���1U�̬�@����J�#bC��LU�Z�Yr)󰡭4��LjQ��������׿����������L���A5CT�����k)$���0��z�ڗd�;\�%�Y&�U5�|�Q�¨LM�"i腽6��袦���^�bqV쁝j8�)tm�#�1��ΤU&�}J���h� LD洞�۰Q�!b�#�c���2_���K�b9��s�i�	��2͡�� �kA�>�ΉS�5���7/�,/v;-��"z��� ӭj�q(*Q��I|hf�'�^"����>�<�ac�����#�����D^Β�p�t[�,����U(`1iL�l����,A�*��N�M��1��G��u�N�w:lg���D�z��b,��S�ҴG����q_�=�T0��.*�i�Eq�h��-Ar��().���j��k2���"��Z��)��LZ�5gff:'/r��S���0s��	#�%�/_~��GO�>���W��٣�,=jG���l�I˒��@�,7���w����$�2�l�2݈I�y��ʒ����5,�nvY��q����H����x��Elԋ�o��W`�`3g�B��Ɉ ���yW��.o=`����^��,.{���~$���6�+l�'�x�)�|���P/H5�*'Q.E�fy����°�:��˧"N^i���|7�xWe �/�s�OmS��O���8����F����P��2��& 䯽v��իP!ءk��͖eS�V��F1Q�p��FtaLu<� ��vb�tb4[-�@e�����_�s,�cǎ��
�PW�~�6I]�i�SPg�x�n������ћ�^k���P,�v�������W��H4r(�MH�  *.S��0
�v��{��^q��I����X���q5|wff�Rc�%�ٙ��o/@�o81$�ɽ�R�a $ɔ���C� ���©����d�:Ne����}R��]MbͶk�2Ͱ��;����W���àS)Za�~�:�p�J���FsE(R=��Da���㟤���q�Y0cM�4z~W�݉�je|���D킟�?�����#J���Ox�� ���ZQJ�`�-��?��3X�\bG�
���,y%D���BT���ۯ�D�l�B9O�jD��3��h��-=�0�,�+x�խ�I�o��E!�(�GU���M��j���	��1��%���/��5�Ч8LdK��N���RQS
�"Re0`z��^A���X�8>#z˒0���}I�v� 8Q6���L��_1P�iV����|#FH"9�HQ݃�m��1�S!�'��tI�⦁���H�L;��u�6ʅb��#�
Q����h��a�s�޸l���}j����b&\eT)W�P}A��S*UV� 1���5��G�\f<ss�;(��2?nB2��?��v�3g��"sssw��e3����U.���Ʀ�
'$=k_����d��>2hg�]M1��s6+ٛ���gF�LƐv'�����J,�xq��)aAF�Զ��Y���=d�����y�(gj
Ɋ6��|�����P��H�3��==���,^� 60˰��[3��W��q�w��VBjn��i��+7�d{�\���\���6&z?R�}[�~��팚�(w�Y����B����+����Ɂ�7M˦m����$�
��̓�����9�T*��kXW��UJ�.�m�� $�.�H�����yD +�
Q��b	z�ܹsXB��t8f��NDrks��e�k;b����mQ1����̏���\��9�XC�����\���Kȗ��1u2,���_��� 7@ȿ�z�wi�\ivz�J�Y�(�K�j�<91M)�Yꩈ[6�V��Ł��}���ò{�����-�}]��]����$�D�L�j�s�HK�-Q��+kK��G/J�=�l)�ݹ�re��8^	�%ұ���� >�M�ɮ�c6�ɢ"�31  �D���^1	B���A�Ls9�P�����)�r���#j�shNB�l_��\wTJ$�H� �#�[�/��(
 Z`�z0?c���i���2�U�Z���i�g��y܇�3Z��W�c9�@
���T���,Y�7�b��tsy�ȱcǎ/U���uL"��F�ү�w&�XF"Z�:&	�A �Z��/�
x�(�Q%F�f�9E���4����#�e�gMPq��E�b����s)�b�w}��a�D�N�"�ޙx/Md$-Mce��
�G�/(�
�Ւ�&�.Sg��������P����s.�{�'��@����fq�X�j�"?H�bCG���Tl�	�At=/͈�juL.f���A��0lr�l��B<������r��`����~�i�!�������%����'�\�>W㋳�_�4�kH뗉�	r����j����G�۪��	�LY��Ku9I:�w�C�	@���Wۃ��7b?�@���^��V�p� ��>V�6�̄�ֲ����Q#~ەZ�R� ��`,�>?y�YxS^H��;��w�޽}�6�S�)����M������J��:�J��5ӸmQ�V[۩H6�r��'I���X�����e4o� �]x�:h1-}�tab�=у�⫯�%׫�Q�����#���4P�-HF�zN��.���.޹�����Vw*�(;�5�$�{	5�îH"��@�ڵk^�<>1�n5��+�r�"�J�lC��X&s���Q��e�"Jdw�,�C��nll���񤐵H��rP�X[[�ʻ)X9Q��s��f�մ�+���8H2�{� (�Q�r)�F�!;qp��-kV�'�+js�wIE8�;;R��TE�̯�Ya�=�1��c��� �pJ�|F^v���ُ˔�⯉�]���߽��t|�ك��F0�PTnNT�R������rՕ嶓�E�����`��׾��K�]] at�'��h(�B*�b�'�����h8)���j��`�a�Q��paw�~>��!��Fu�	�E񖐍��^������P%|lĂ��L(�%X�`�T�8y����- ��q�8
-`����wwl�A'�=#�ˎl/G�*i�qCs|-�`꓇����0(�~�V�|�.��k�Y�/��).�FI`FjR5�k���~��qd��9�B9���gόOzW� F@�Q�$�&!�R�e���S� ۅ]��u��	;9��"0�>��9nG��pK��ж=��sZ,�B0��B_7�6EB��7�O�@%�#��EVFav�$ �p<7�g(,�i���?lf�8�?�+��0�L��r���Aα�
u3��Y��'�ɫ�c (�C1nS\�aAW�q��d3��+� ��`L[��@��P�!SK}۰}1�T�qh��ֻTq�A�+c��7�X"�$�I���-^���Ӎ���M�,��݁1L�ĪA掃��B<vl�a�-f�
(�J(���94|���+"mB��e:nͭ���+��r���Gy�s~~��9N�%�v��o���{��$���V�?���%l;n{����e��}y��n*�S\�Yɼn��md��N|2/r��sѯ��dtk�|��H�^eV��	G*&9����
㽑Q�sI	_�O���[|)�|y���F<���g9�P6��d�9q�+���"f~<ٯv@Er���� �>�i��J���ˋhC$�*����+'B�����PQ��a�y/������8�~ԙe{����q��Mqȴ�hp�"�M�&ؤ<���<xn}}}ii��lY���5F���G'��ԟ 2�wD�բ@:fF*��ݻ+��,��$i���M�s<[.7�Z{��\j\�[��v*EE���.�?���J0*�P��j��|���4�d�yxU�r5^$Q=Tp����i< ��8e�]�~���Fxa�����K�,�I��u/_����?^���ła9P:��9�(r)�V����M��+[��}����;�p�<y��OhE+Ұ�CۈuR��������Չ)(.�SSo\�|��w�:0;�������{]t�wXJ闑��2�fw�,nt���vz	�?#�WWW��S0�Y8��;�`6]%��R�V�b�}O<�Z[i���a��,3g�FI$"Q�5��
������70R��K��-����pj?&�D�����q�&��8�Hв�t�ݓx4N�r��ܳPU���D�]��WUH#?W�A݄�= �(+�D���+��J�6�y9L(e1Q�609�]8�b�:q�R74��SO?{���v�;��/�ؐ�N'�G ��\�*�cXA>5$�Mv�I�7�8瘮�fe�����7b[�
�X��S"r9\@�w
�N�R�B��B��&W�'Ģ]�7;͎!�8ĳ�׈��X�u5��2��2���9��M��#�D�6��lWvDZ���$��Ң� w3���JH1�!!<rf�)6)G/���V���~/��(�"k)�֢�Yˌi�4� �l�TK�i�z�:�f Xe �ia��Lxg
2���Fltqwn_�M��6��q�iT�)$��um��"��s����
T]D�l"��)=�L�Z������� I���4��E|��ͦ��S'���肝F�.�)��ȌV���y�q3�CQ��ۉ�/M�VaRpX��(
)��B�Xc��Q��-�X�af�0���s��,6�`����Df�������n|p@+0��������ϳZ���իW��=�O���X~�c� D�8��gmm�#?��a7�r6��l}���Jj��/������H�#��m��lSSS8ƥJ����"M��B�%�W��{�{ײG�{��L�?��SԀŜ���R��šv�3p�IԔ�;8�/�3��8�"�+��%��۩�x��ǆ/W򰁂�K�7bg3�ȍ7� ������=ccc�<d`d�)a �M�r�V.8Y84G�ʰm0����l��\*��$R�g�+����d؄)�p2g���s0��=��cf�G_�(8*��|y	W���<� ���%lR=!b�dPZ�+4�z�Ԫ�����@�F�) I�D�=}Gh�N7�E6��F=����p1�N޿mJ�xxH�̵���C(I3�M�C볘��uUH/�aye9/]y&�5�j��;�dEbi�s2O����Kѷ�,}��T��C�L�¹n�E�n��I�aH���Z�~��]����:��c��ѿ��yꩧn߹��$�.Hb�7N')M���$�T���W`�O��ʯH��s-\':��P�q�si���4DY?�\cfHn�=�3m���8=u���;����S�N�M������ql_�u���6�q�[���}hA�@haa!#����*�a�
W�L�W�j��`�����톀H>�p�ZI,���H
2j����P	@��Iǰx<Mf����&R��N"��]Ƞ$�`�YI�Y�ϫ�c=���0�ƫ�����S��"JdJ���m��Ԅ_5�n�$l�1M�C!a���+�x��"i��;����tj�Eg����>q���4�r��IQZ��>L�8��v�?��=���Q̼W��c��w�����C�H�bQF I�ĖmR�+,�c�kS��{,"/>�h?�~/d"�D�l�]-��\ˆHE�����0�a�%�5iiFhAQB漒i,�;�#G��sŜW�y>۔d		�3ټ� %;�`��*x �"s+�@̌⾰�lӰ�ur�(�N�{��+��z俙x�F���@����`PW�0��縘
�ݎ��}�*� E�Q':��n1T�C!#@�<^'�������yb[����ST'cv�5��(��q�!Ssӄ+�d��.��DV��᱃(0��+V�����7y���eR��Lwl0:%ӳ����J2�P�4+e�D#DYC�� ��ڞ�����-���������&��q��)r#Q�j	�B[����>z��1|,����sXVH+��}`��_�"|�M���p��!w?���o6�$Y�j��/b��f�4[el��uv��J�����mf�㦖��������f�΀��?���bx_�u�xB��:��V	�����G~Y�˖�,�"��N�Y�I�������.//�A�E\�&Ǭ�
���i��#|q��Sj�.�GX9���/�/|��G�(hgS���y�Fx�r�.y�J�U�� �!�P�n��Q�K��I�a��+��	���2j�.�.���Ln:�t�
p[���|�Yn4��^�Tw��P�:qk��mZ�S����z��a�]� S�8/'��J9��j�\������z���;w����+�')�j��$C�EE��kׯ_�C�Z�̙�*i$LG4<Θe%Q���|�4<q���<��II�")��*d��J�P��\���x��"�ɖU��dϐO��ã�/�^��
��Y� ����e�e���5���D�Xg\���tQU'����nB���s�=�����~�G~xf��F}���+Q���k�NqЩĚ��s)�A��8֘�زە���&K�ry�@��_�7?N�6YYY1��9�����=�,M��/��o�8yfg�.��. "sE��	Q�i�l�.
�TU�����-�J�Kt�J�_�"�Y�IQ��%��v�q�N�I=��훿���t������.8��}�����9�	���j2r�dav<1�$?��3��tc�B�Fuߖ���^��R�ٯcT�m����-O$���a;|�Y�B�rxBH�:p��T�E���=zg1ã=�fǍP��}��a�����I�~���|�87�w���mZ��c�9���]*�BQ[bh��8�bM6Ua��p�I��J Z��Ѱ��"�G/	� O��\wl�H��v�U�H V�Ȳ�(��x'I}�2�h,Df�-���Z�/�R2@D�LB�� -Է�q%�%�D�`5�� ���I�oki��J�%���t����[�"������ꂋ:�#ʔ;pR
{O�������h�X���Ѡ���E�0�u7bS���2J���f ��@P��Ѧ�2y��H��FX�0�4zV�(�*��S%�>�����ih�;[!;s]�$"-ߧ���u�f@J�3�)�X`*&$N�J�B%@0E��D�fٺvJ���h�m��YJid�ٶ߮��J&�PB@��vkWx�Q<+""ĕ^활�h�:��QP+�ڙ�5��~F�H�� !C;�a��%H� ۄ�H���!���âAΪ�ܝp�j�G�����ex�RF%5�50�xƐ!��,�pL'��l	�:&Ͷl~FU�z�?6(�-b������?�z��{}�v��n����k��k����c%I3�+�rO�I̐��Z�������`��>}z~~��>���a%�_|��7��	%�9�!��ج'V�d������/���))��A�Wc&V&��T�z�d�?�pKrV��m$�����F�do���?��?��K/A�Q3�^���쉶����0:1�X�;w�0�2F��������Cئ�5��^[[[����u�y�>�,�8����nܸ�Y:z��I���@��D�-��`5q���A��®`���ĉ�o^�u���N,ڑ���Y23S4m{?8STLŔ!Io8���K�*5��f��l�0ms����5��a��QU�c� Hw1G��@��9k�w�c�e���4��i]|eޥ����?�F^�R|�;Ւ��}�7~�7Μ9�����*W*�(��+P�f�Ȓ}��^	.��10Z�\�t}1x��?�w��ۤ\��|��!d$��0���@zs]��J�7�H��Nf�)���)v��)�;5�����N�:,��o��M���~�/,��N8kǏ�����¤m�P(G�xdm�Ht�!�\���[r>�,�J6;�VA.�>���6�X|K�5kn~��g���!n��n8���,�6�F�(ظp���N��-Y԰"���$d��%���b+�M�uz������*�c(^��2z�x���H̚a�T4�z��f�Z)���s����0�c��(k�\�ރ�������z�R(���vi�d7����w�="n� U�K�y�����ælĝy8���w?/�$}l�nx��	[= �,�;�Qyte�=�~���4C]5cl��La#�T��o����V �U���PN?�x���:�y�L �i�!q2G^+��?L�����������3��,OD$!��%yD2��)9�������ɞ��pK�[v 
���D�,�Rf%�|�u��n�nݽ����,j_4�(
ܩ�H$7e�[���^�eٚc�qo�t���nW�����f\+��70��SB��>'�K�|���R��䐭A�!���̳@�-*��r8	�m�������D�F�*x.���E�!X�I�F�ߙ��p%��=<�i�!�r�?ӄ����ȡR�LD�4�����iE��C�#/�]��Z����hRP����lf��*6F	��門"���1�"`Q�Y�FӮ��b���cM1a��u1�M��#������J%4X��Q����g�޼��~�����X���ppRUY�b�7)�/kwZ�^����$�z�����nٶ����dq
C����k���;@1�%��C��:;�����_��_�W�;�e��`H��V�&40�qpd�G�������I|cc���[9h��6I�*��9i����p8���L?`/ݏ-�eK��叴i��#]�Z-��)&bq��X�n95��|�h�R`��qN�7��x��շ�~�8�r��5�$&������c�a��\����'�b>EH���'>�	�&^D|+{���/}�K0a��R�pr���ۗ.]����z
K	��'����jĨ���W�wb�qA�2��|��w� �pS|��~��p�����!A���H�KF�+3��x��h�"����*�x����#���@l�s��>\�����-'y�� ��`uVVV ud�?�g>�O}�S�xa����_�|W���g��ߎSy�2.�]&��+�Z}r�k*j:;;;335.��A�
�b�sW�6M�}"2��@j"��Q��R�>˄L$ᶸ8���뉌 ��t�Zmvf~cc���,A4�������Y�s�a~"v��dO���n?+�����"��Ew�ፄ;Ba�T��6̏������X��z�9s��=��֭[���u,�0�|Rp6�U������#���򄞔�]9Of��"5�WU��%s��9�vw{�+��gj�iò�\����k%S-�x��:��\+��pV�N�ˁ�Hd��	��,��(aO�)�t-��Ru/45���YD�ƌ����Y��<�*PӉ8W����ye�f@��XBam��-�k*]�9J��/����H
�OI�?b����.j��R������~��#'���*�C�?:�uF�~��PZ	�!��I�E�0�$#�#F@q�?ބ�]h�wPo��X%�B�-2�B���D�x۷Q13e��V��ۡ�=:�|�g?9֜���9Gӎ��j�XƆ�N�
�t|���jgf��p0ܸp����Hɭ�o��_��:�d2�3����0�����w�.߼3;>^�s����gN������$Yɭ����.�z��͇��7��ʱ#Ӎڸ��*���
�>R�rS�ېn�p)�R�~����Z��?$*tЙS�{����:�\�eQ�ᯄ&VX�Y�V�S����޴�Y�D�j�M�L�(�N�
c�@`��.�l55���v�7k���S��ɹ3g����y�e�����K�S�A�7��X�u��ѣ�a{~R��[6l����7	�Y��/��Vn�j��.Ζ��\�Z���i֚�'y7�/�c���fQ�T������7/�)�\��r]�r�TU*�}	��J�Nك�6W�^����T�Z�91Ѭ�TO��3�I� ��HDf1>�ky��S�Jd|P<I��i�|�c��Qu곡�~M�V���?���۵+��Z�Y�V����J��Q�7m��܊�o`��㨽^�>Z*Gq�������~�8���cc�OaL�5��yQ<"��MV�K3���ON`����q��'O��ad�'��j�|�ט�Q��zbb�������!{�����KQ��7k��=ߜ��f�5��z�o��=�G)��!��^L���j�۲R孷�b�y��}X��{0c�%�Ň�t��L>l\<���KN-���W|�ɾv\�
W~��9���R���ѣ�60��ܹ��@����G�Wp��ş�� i��<bG�.0��1��d�?n�##��;�FH#8p�`�4����=����f�5�:}�@�uEB&��s���4�$����/�g�O"s�8�#3��E,.�m�3�j�r�".����������+�30���o|�o0�|���\�%��$�H��>6��?����_�]|�������j4j�r4ʉ�t{}�>����V�PR�ޠ�+ҲĢp���'K%J�sݲ裕 ��گ��k[��_��o���.��;��ؗ�b<�xI;�>Ǆ�!|dmL���{s�����)m�'�ÿ|�9��y�1���LJ&�K1��B����z
(�5�,R8�KN&0S�S
�!�Gz4"�1t�;��7��M���X�~��{a���Tp]fv�I$�H�u3Sf	�'�����t�-�P������{� �9���sn�W%���-����#�&E����m)=(�bUh1l�/G6�"}�������N���S�J�Dqe���Ʒ��w�,�tQ�)�ɄX2
������I1���ӒW�}����GT��<a��a�u�?��1K?�Gr�IeP��L�e�B���d�$�J�ԅK6�i���=B�s8�&"B��\��Ɇ����j�J�B�j�v�E0�u��3iBF-NQ���r��kaw}�Y{��qS���'��%�l�1e�Bz��I��"%ݭT�0V*���~i��K��a?Y]�9v����B�V��Z�"(Y��:�����Z��cc���'v5�ʉa�k��GftMu\�֧��e �x�;���V͍��׿������/6���1euj=F�O�؞8�u� �P����5h���x�����YMuk�^]�����èR)AB�U��N(NP�%�5to.�7�������j�ߋ�z���b���9�0�C�w76����X��K_��fǋ�֨���2�_H���\�fj:��X��Nk�����?����4�����cGOM�N���c;�`B+�D(����7�}��c���^����;{�D�6&�R�fR>RR� 
#*�����ܾ}%I����%�<	Fl��"H�
Y�R0*M�̿y��oa~��ÿ�ꇸ���X�R��h8�4OU��dS�l����=r��E�"�w<r�87Ud:��LC�I��0��j���~�?�������ڭV*�i8���m��|r6CK��0�a�b�JH���
��`�o[����d��Sd�n�٤xi�Cֳ�"@��]A�(��ǋ��G�M�.C΋XZZz�g0H�3ҕ++|x���Fζ�2����K,Fص�I2?F���Tl��z?`G�����H@(�L��v�L摯���ŦƥK�p�~�~k�ꫯ�0�>��Ob�`7H;�2,�cǎAN��{����`��T"8*8��
�b�$��s�=��7�Il'n�A�T[[�ϟ�`��92??/��0&ćq_|�1�����v}�؆ÿ�z���0��"�E���a�*��t�\ŶHEv鑭�C!�H�I$0r�g�{�|�?ܘK�.q�tP���j�Y�V���
_��W�g������ÿ���ș�<�����~���v�������6g���e��t߹�9�[��&�n���S��q���5���z���ڿ�7�fe徚�\�D$��8���g��ٗ^�����%��0�VZXe캵�ͽVG���RE�\瑈��� �4�o��GQ��b��<�߿���d���pP��R&\VEC���� Ib�8,����?as2YGۊ=j?|ָ2�'N?~Cz���WVV���3�rKJ�E�n|��P!��������sh%� ���>=��$x����#Ll�f�iUKnF����^;K�tФ���z$�:x�J B�5�}����1"Y&�,��U��)��ݴ���c�E+nɑ �]	t�:�[���� �茔v�j�D�]f+�DLT�z�0�b��2��G��p
>���mm��{�MQH�>Z1�$#B��a}d.o���GW�Ӡ���#Y\{��D:�if���vc�"y���YJ����#pS�g�̦(���Z���R�sve��<_��e�,���Y����|x$��1��2ɻ�����0YR��7o�t+�����VFݱ�Y�K����ֳ�#����z��{E�������Q��խ���--�]��A���J%�[�V�\[�︺e+x���GN7�v��6ַ=?k։U�����M6��LZ�7n\[lTf�ycf�6nl���[f�Qӵ�{{�m�)�S��ò�����qT	��ԩ㏝=��ej���A�$�GİD�47��U�=�0��S�O<{z��W/�X���ƍ��r�91���'!Es�D�;�(Jʓ����Ɲ0iU���k�A��ƌXAMXњ(�!{4K��\�t���Kg��=q�hɴե{0��oH���0�]s8�@�����W�UjUC'Z�"�Y-ې{���þJud�b$T]M��j�ҘI貝������k�kF�����e�޻�������P8��mY��qB��n9��� ���Jp���jkW��X.T�.��Ie�8����[7n^����'��s���՝� f����5,|U��?"BB-���W��Ͷ�%'��$�)����]���Q�TN}Jn�0���v*z����b,n�Z8q�:�:Ԅ�Ij��[_�qY�#��J�r�٘\[[�k����y���~�I���0�16����ac|2��m�:vl��l��qL��ЁL�n��Щ,v�w��б�_�W؎�-._�3�CIAƂ�4΂c~9�%\���m�J��&�+�I��$�q���>�="�d�����1�)S8��ǉI�a��X�O?��-^ !<N�#>��1�y饗`�r�=�
Qg6��䩩��xݽ{��¦�g?�YfR��.�(��s����Eď.\��a���"��0=1l�C�n�+@bco`�����W0=�G�
&|����D)��x���s���+YM^�zD�Y��o��Bzaa3�60�Ћ��#�w��y�E}���	����}����g��$L;�7�|���N��5�]q�?��?ƿ'F"Cx����.~�i��7��|�65�~�Q�WA�mԚ͕�՛7�//ߣ�"���iu�(v���'�10��i����	� �H�T�f��;w�w~�w�Z] ���	��w[[�>|�������i�L���DJ~@k�~@<�׿�u�v&s�0���KlU��x
�v���N8����J#I1?��	S�!-//s�1Ɖ��EaL�{����� ���NHk2�b
�.m�ZWPA��r���s����E�&L�{�r !�^&����
V��b�R
aX�2���֩��.�u�p��K�yle�f1C�7�aX"�m_�k����ع�h~rm��p� Ke��<�B�UӶ(�.�/�q&��x
�F6M|^�Ɗ���Z�έ�/�>?���@b�A`Av��m=`>Yd&�&�:^� ���r�7r<(WY�%+)���	��U*�.��K�YX�1;礢�,����.>ؼ,:y[p�2����z@�k�`�8vݱPfa*h!�a(XX���iW��3��.ʄh��G�;I��]�xx�b�pM��Q�-xONn��j^�U���J����Ogf�Iٙ�v��=�G�O��k;��{+�+~�����n癧�4k�o�Uh��ף82�T]�ֹw��?�g*���k�kC&z�ž(`*���i�WtT2��|�
K,{,ɴ�\:�TvV�Yx���,�Q�;�@�=آ	eĥ~U��n&�7�W�瞝;�΅����^��l���޾mh�u i]�r"��$&_�F�x?mVk�	�U����MU��j��8����b(���Q϶�t
2*O�H�-ӨXz���c�������ݽ��v���z�i�C�W��^H�dY��q�&��+�	C�*[� ˏ?6ulfr��M�^|�c_$��3W�����V����4�~��S���{W��Z������{ׂ���<�ھ���<��9�"?0m7�U�\�����'��::{���cˆ����F�	�^��V)�]�oOq��O=�r������f'tb%�����p��@n�O���ƞv������EY�5�'ϾXV����u�TS��2�(�	U;DzS%Z9|#�^z�������Z���+�������^8�S �8����F�`��H늨�dc���3�x�Vs�ȩ�Nb��ӭ��+NC%���������uo^����`��y�v����2�q�1�dJ�b����tY�p[��ɦ�N}
rLU��n�319��Y`R+��hлr�M��L6��C3��_��>_o��pY��+Uȑ�j�W�76ַ`]��J��h����i��%�_��î����|e��S�/�U����6�hě�[\8�P2�)�~�nO,'�ܥ�%�=���󄽃x���+S�Q����yTX�R�}�ˆȢً�3�3�����V���bX��Y��S����m+�"a�H�p��li��:%����B&�33S��<�03y�r�v���p�S�����2'G�t��X��a��A���Ef��n��)�x��IL����>����c0�8Lύ-�U`��N@�3��'`��]�.0� ��ln�Jv�R'j6�S��A;�Y�w;{Lg��D�T�HJ����\ǲ�♘N�UtKD��g�rDA���=Ԝ��0?P4��-���Ѿ4!d�T*�V.Uf�o_��ؑ٩�����C����9A�&Qm1]%�R�v�'5u͡7�E�U�5*��-j'�N�<]u���n�{�w�N�}���S�zUW�`rrZw��%����v��"�1ݱz�G��T�)/��(��-W�0s�~{�46ט�7��ڌ�ۡ�O�eٹ�����?����+o�q�_����n�UE㔳f�h*u�����`XO������ӏg
%���8��qxU��D��f��<b90\Ⴭ�t��N�4*P
�^e�����6� Dd�!���B�C[���诊�/2�`kkkH�=���qЏC^�TW�g	�6��*	���UM�h ��,�hzE��']���3[�<�Ra��!%7dZ�&��ps��:5ǲ��ʈ���U2b�^�z�t�;�ebi���O������{;a��7-R�!L*�5� M�$"��D�nj�*$H��8x�Nt��(�c��j�����i�,p�D�z�}���-��(_��"^!#3��[��Z�
}��;{����ką���U��5ezuc5<��h���;Ö��
�����O��O��+�f���$\�m�#2q��(K�Ñ�x04���b�b
���=a��;�>J�*�<E�R�%�#W����Y>_YJB��if���A$�����VQx��b�Z��)��%ĲvP&$
�\�D�#zb�
Ie9�k:EK�Ft�(�"�U���� mC{ݘ}��Sg`g�-ݺ�t�S=����,�$�	["��\�bL���ٹ�#sGuU������u"�6�v:~���j�V2U���LKM�ʩq�c-�7�Ju����R�~�NN�ǂ�P3-�(�#ՠNB%���LI��8�d�(�-߽���:T�qza[,//���D4D��Q�����t'�k���g�&�����:�ް^s6�R�M�y�p9��2칹����k7n\�vm���'A�������R�'�*Ո֣9�^�M@n���G'�~&;������e��tT%�ZS�����p�x��]=jo޻{ou}{7I�L�����{o���n}O���JI��dj��O}�rezan|rlzf�6-���Xu�:U�J�{��Ér]�(a�z~����騤o�ٽ~�2FS�N@����k7!���Q_�l�^��a�\��9u���<nT*;�SMVt�[V+�i�Yr-WWL� T#��Z�U��z���|�Z��|�i��7:�!�SK7��i�E�X������N~�N�V�N��v[;�{~���A��XuJ/��ԫn����w�-2�b�%����n]�zuS;׌0��f9�-}�����?zl~|���ձf}an���3�[e]�ۈ�ܙ�0d��b����W�-��S��V��h��O����̱1�j�.�ņL��uj*Kd{&I"E�=�����������7�!-�w�EF���6���"�z؎\i�?�"�`Ξ=�s?�sł񽶶q�Νrٝ��406:%M0˷J��0`�"�$ۣ�����Թˊ��f�_�J6�,���	�d9ƌY�3�� ;��nN�OLNC�rw�ag9�7s�]�YU�k�ƱSN%�D1띤�~Mn��b�#�r�עpd���y�8�B�:9�Ĳv�T�����ꊾ���K9r뾱��ɜ)��!t�!;���*���swy�c��GU��2���A:FaK�� ��;w.�iip��N.;��������$��JKI��O��Ül����1�{KMT��3��x�^���e�����Շ؎mWba�q�S���e'f�P@���,3b�#����SO<~f�^wr=��,�5��$`���/}��?�����#Jգ�$�!�H��dX)���۵Z��p2a�g^-�b���x��7޸x�"���{�,
��%�-N� ר 1�e-��7���2���Y���̮s�X�Qq�Ē�|�4����'EDĈ`CY���kznv���q	X�~u;�$�g��H��������x	�(��S(7�9DN��1U���rC��]��H�R�0.����Kg] Ӷ%
����9CUI�/1�]�Y����e~�<��O���%l���ď44]C�E�f�5]�X0:���U��YZZ�p����
�(�>��1-C^��	ݻw����Ͽ���I�vʞE6FyZ�O���:H�H�Çku=���p_��Qf��w֨�x6�):ȕ��e��A1�>K���=�\:e 
k��������̳A�|@�4W3U�jm2���N�)e.YT�N4י�Է�}��P��}���WWn�|��ϼ��r��ǩa�\$i.��<պ�T�SR��}�����]Oӭ(�c��nւABg$��k��2��~��)���^�6�eJ��^����|�<>���$�i�9�y�,��(PR�>�TR���{��-��lw��ѬM��k�����`
�U��5�d؉ݷk3X�Z����7��|�^���c����~n'����luL]q��7���o��+B����s��k~�g�J�g����,틱�;a����v�!�4UKb�ųͲ`�S��`�c�sJܻr���-S����%W3��݁�i;�\�ۑS*� �@Й�V�V��-�I?���`o�:�b۽~ �t+�0�&!Օ����w���,,�Mχ�>T_�^���;��X7,�P���P�������U���f�v0P���>�j�mP_ C���1��Y�zdhI0h�6��^�R��!4�N�����4��8��R2j�(&n% ���@��Xy�lo�����v�c�sNm+'H��1�Y�p�ں긊O�j@d*�򨈷��{+�L�� I�:�"�*���L��7f*�T�Q��ݲ�@��J����&������ٹi�̼h���K�jmrv.z���V����������
�� @濰g�;AƖ�՛��gO?~tvfr�^
��mj튉��vl�0b)$�js�5!��`��߿ϥ�?��f�	�����W~4�ʿ��׮ݘ����k��B�H�<v5̲�q�>x�
�@h��ͣG��:�V��������������9�������ˍ	�Sc���~����8}�ZkȢ����H��K̏��������rdzI�hY�-�e�Df��lRĩ8�iLZ.���3G�D����p������y�F��l��j����M&<�� ��X�r�+'����]9}3���o�:������>�d�`��2$��ϔ�<Rj�L��-���#C�>���}�S�����}���񩏒�Rͼ�$W�w׏��#?c�c�ԁqu�G�#U�뾥�LN��,VՊ�$K�[7o�����֟c�a�b�f��Z;�%N�uo�/iʱc�l�� i��TC��p�% ���,�o~�@�gϞ�Q��s"�0?I�e����������D|h�K#��E:�:����p69����H����(eN�o�My5��Ği(O=����<U�5�]u54��Ay��s.��'Djiz�+İ��X0|\��ƌ:��ݩ`ʾ{�y.��y����2�yUi����ɣWd�QŎ��]��yR�D�vc���~����I$D�ۙ�)��an�B���&1Wa=�r�S+.T+U*���ա�����ݻw��tsss�7贻#�j�Ģ��0�&�d��Ll�a�b]f�NR�WAއ��#���!z��7#������>�a����_�?�2�;���kE�(�6jB� ����,e�
�_�{^���R.*N�r��):���3W��9� l�R�	#ϴ���f���_<���?���WE>x�QaLkDg�_��0���[�|�[���0��H���0��� �\!�f�֔:GR�q6j��`H5�1;G\�|�{'�>�/|^���`jZ�u��=��
y�*I�|���o�;��If�z�$��A�VZ�}�jUL�k��$���#��0�''4�Ƶ�V���3���j�+�U2m�ehľO������x���&Q�B:AT��X����6�(6�K��L�8J� 	c�p��u;�2<3�wj��G�]~�#/P5#�M�G���"��P5���ƕ+W;���OO2��� 6l���C��҄%W���`8qZ�8Coa�5��[k��]�=vvl�`�b8 O��P��E�r>�J8��w�nc�G��0˵n��V�5k���ȋ�<
�/�,!pɺ���#7�{����R����5�V{��)L]�r{
���5���I�^��+Qs�nkk�.
��N7ו�Tcja���V��s,{��´���S�Z��j�� l�v&�>2;9����'N��'��we���N�Z�ǚ�VD�m��N{��L�~=
2�j�Rn��C�M�
b����W(�2$p�Aj8�c��*��ݣ�`�Ҁ
m]�0�Թ:3U�R�r�� ��o���Y��Yv�;���ޮ��o���N��DUN��"�,%���W�x5��'_�0���&'G��	k�L-NE��Q
F�I���}4�qgg�=W?r*�sğ������<~�8kz\|~~��_ru
[ ܷ[�q/�:@�̭�s�<ikkkDaT*Ɍ)N���^��QΝ;�u��yF?(�@V�\ս���naa�ĉ�F�\�q�<0�6�cqp�yDH�)�a'MLLpBz��͌�������^Un(��8��)��r�ť%�n֪���ɓ'{�ޭ[��y��jL6E��GA2px�Zd��$��vW��&K���Ⱦyޘ{W��3���/c�cCJ�Di3�o!J�>z����~�fݠf
��}�D"@��[�Gf�)ѬWr�������ُ�@Ľ��*uW�I�p�#���H`��� .O%���		-ײ���o}��0�z�*Ŵ�1�r}�"b��%3�$�����'�C+�'��p�~KiC�0��w���^{��[&��4�"�T�C�H��D�Ke�B��B�u!��o�>�������ċ��<z�]*�Q15�}�/�O ��7^�~�S/�����?�1�)Gݡ��Xj���FA,p��8Q[�2)	�dH��(9[�n�
jɵ��	�vC*
�E�'��S�0 �4YlK3�A,�D�O'	oF�^v@s�R$=���t&��%E��;��ѫ�D3���7'4������1x�r2�r�s9�z?�*ƽ Z��` -�>8���cv;ݢ�?<�+S�;G�UN�� 2lz���8�GT�l>�6#l6#y�ũ)RQ?������<�9����<�v�
669�4J+�Dv~&c�"��0��(J$�1�/�:L伾tL`�4iu������(������5y��|XK�������'��}�w����;2;}�8Ĭe�yj�뺦�~���ν;w����޸~���Nɽvw�!e0$�Ha �	�H�����JBi`T_!�&J�YZ�uj%wog��[��j��cG���ӝ(�C�4UW�H�:���x���o�Yv�R������a���ǝ���aʪ�{G�<`�*�����k�R���n�W�������O����1uf�嚹�Gl�7�x�¥��f�9c����:�I��?��� R;�G!T"��Y
�V������z�\�TJk��������Ԃ�:��#�G�Q��2��0�����o߽u�j�0��V�3o�{��l+rZF���^�G�p��{!f^Ӭ��ؽ4z���*�ӟ~�K���@zx���m������g����u��׶w�t���`����sJ�*|�Ea�Z pԏ@Sm�^	� �9	�H��hss=|����O�͞��<���vGѬ��yx]-�SO�޸�r{�����Q�yYc3��0�[��0B�CW�σ5����cME� �a,LN�ݽ}�տ���ѩ';z����˛�F	�ް�J�f&�}�.]�z�"`������2�X��ǹG�D#�
C3TDN���9S(��9w77.]��B?���R�N���!�%d����z��C��J��!��PW�F������B ߈z�)�XO	�!�=�i�A��~��ʤw���\�DjR!F
��g�!e&ԉ���k����2h��F�q��1�*ɮt�����	�	&��p�hbY����v�F� -..�P-O�	�q��g�>�䓗/_�!)?M/�� �+���U���}y�^��J]�%KӜ�E�,��X���MõU�L�ȭ�
�}�#�I_\N]�������1�C�z���7���>���<���4�f@�4��q�'�U�L1��֜�Ħa��*ϳ�T#���a˨��NNN�9s��*�ϔ��!9�Ɖ�𜼟���&e
5���[�sv������+W.][�yg�6���'�k�1��gʹt��پ��"����Y�}�в��A5Im�1m%�(������z�|^���nwv�p9QEN�r��,�`���c1��F9dҰ�ʃ�9�<v����oooC�2'�K!�����`�R��
P��G����M��q�Gx��Gn9���K�l��x�7��#�#m]��-c-UTʵ<K������������n�;����P�@�4�dr�3�&j��"L:{�8�g�y�y�6t�4V�
�Q���zlO�U�,�H��LMM��R��bW���;�S)Ś�Գ���dJBq!�y�����nq�I�Z�FY?Y���m��������+�+��۩�>�2�����!��Y�|�S2.��A8��m�
���ɱ_�p�����!c�!c�E���>�����?��SyP��"4ztݭDS��)ߏpD"�b��b��(��(���]֡I����DY��h��@�8�5�<�A�B,^&�ZTr�橾�O&t���Cѡ\���r�Qv�%�y�S����?�_����寜={�����ЩŃ���.�}��ͥ�wM�5��j�M� 
| ~��G����!ezn�[�SC1
Ui�!��%_)������?;q�ԓ�~ĭ9����f���{�ݭ���W����ۆV�a@'jwH�{Ȇ��nJ]!o>�'s^�A� ��1�<����T�n��w�7Z����<��Po:&�vtá��A�{�����^za�>N�bA#���G��ޯ���ĿxH���� ğ���Jٽ��w����~���ss�rZӴrFQd^���[��ߺ���4N&��vv[���;I=�7��X�nA�&��e���@�m��B��|_�ͳ�?6�h�'(�2���KC����Z����o~��:�Tw�ݶ�-��nH"�=�������f�ե�'��ٶ��T\I�Jz�ֽ�^��S�Fc�NG�R�۹o�yբ���Z�����Wo�[ԚV)�M6�y��{ �(K�׎j�1�PfL�*
S�$�jꎊ)s,�+�ݟ����Ш���a���Fk�����u�|ϟ?�{�ؑ������8�<c�Z�HtQ2�]ɠ�����]����'�"o/��`�5��<c+�poӰ\�2�U�{A�w=H�v�^o6jM/)9!��O�DO]ڗ��Ŧ%�v�H`1��2,�.5�M]_�D2�g�i�q�C�"ꆌ0s�8������G?��������r����y뭷p���if�>}�t��S�ǅ����o���a���������w����/~��[�<}mm
����,�\A����aܲnu��&�]�Z����&���I4q��x��Ǚ��3�eT�����^R)H>�A��㸖]VR�G6Y��h@��]�C�
Dר�I��p3D�=��g^���?��GO�S>�ybĈ)���l#�d��p-p_��Қ3�Fc�[tzz�z:j�Y���<�:����9���"Vr�,�A��n{wk~~~�ȉ��y�N�g:��V|?�6��6���0��(�+vw2#��%����������Ǆ�T�t6�߽���BJ���aw:�0Hl�%f�vW}k�؁U	:�>zye���mʟ�8E�3)�Ó�Xhbb��{��' 1$����M�1gx6yGҥ��/.%o{�#�^-�{�-�C.�(���rL� ��ԗ-�dA<��aXk��Bd Q
�?�y�봌�x�?t��faЉ���e3s�l>�7n^[�X~��W?��Ͻ��K�F�J������2� �X&{U0~�#$�����N���L�f�}���@O�D����o�K}�H[J���H�=a����Z�:Q��a��o��������~����c�fg�1+1�1�)�J\�"����L��;;;��(3Qά����%K�x��^��Б�ۈ�b�<L|�¦j��n�|�����~Ż�t�+���l��AP��O10%�=e��b!������ ��M ����E��v�'��_Uz��u.�¾���} �^���O����� #�}yR�O;�`�CI"��3,���jGg�~��s���ѿ�Mp��Jɵ���dwwmee�⥫�;]���Ze�;�,����
|�i�oي������G.t�	~b2�0RҬRr�(��\��n�����.L�_'lo���Z�����v��l�T����T��YJS�)8+�t
�ɋ�Gy��E��E��T*Z2��������݆y}���W;�����{W���v˥�i����d���6�}`z+	lt~D�I�'�賱)!3UIt׭B�����7�<�������\1��:�wڻ;��^g���r�֨O����AIR�X=-��[j]�k[�MĖ��U�/	��[]�[���Ͻ�k�w����<��%�d�������s�.]������af�E�l0�U`-#�|!Y6=u<���҄"�I�U�ja�ۖY)�;��w/n���2��ϔm3��N�{�au�ݛKw�__Z_��ƨ6k@v�F�©�=/�Ev26�ip��}�C�V�8$��(�M��ݽ6��/�����qv~N�\�Q��o]}�r{�<���C�,uoP��Bo�2�u p��ڎ��i@�癬�#߭��fq�מ�����{�o|�����_�L�O �����K)����q{i���6�j��-̏]�`cS�J3���pԅ��jg���H���J�hʌ��3y&#I���~�LI���eV�L�N6e����6ê���7o����s�~�wwi�3�b� @��+���,,4t'����]6�pr��~���E��Wx؝��G?��������5,xn���?� FDZ��ٳ������/ݹ��/�|��|�%���jlI�'cA�)��W+ź�^�ː��ə��M�����>�Z�`���|V?z^܏����X�~�O_��+=��)I#�U�%F*r)�Ӳp��6�����jZ��1 
��s)]�s�qƗ��±-�	��Dc�YX\��������ɓ'�����w�}���{������n7vJ�J�4>V�S{ii	`�7UN�ͦ��"cD�4�iV��À<O+˷W�ݺy��ҕٙ�'���Z��o�{��77w����2VB	���?E�م^\�1]��G�$o8,�7&bv~�p+��I߷tC� e�n����0��	!G9T~"�uaD��;��p�������B׺{-��0�Re­Y�؀�Z(��fi�R!�j����3���<��t'Oҗ���W;��Bơ�lL3��q�̳�����ś7od�R)(�6zL\��,Y,�8r \�5b��	:.�Г,}�0l&�~
~>���X�1>V����N���{�.跞~⤦��f����.�fx�0��x���b�q-Є���J��F����d�m$z8"dvX�#�<#�*�"~("�]�wX=�p3)Vv��"�b�^�s�4�	}zz�^�ů|y|���~PZ��=��}�B����� 	nb�����_{��ϟ�\߄��Q2@iF����*��0����yZnT�u 'X�33ث���{��`���s�Z�\2���dSf6�uM�e�řjP��jf������s̙n�:�t�@@�C�S�\�3�4� U��F#��}}fv|�^#�-MZ��0�U��襧�~fek#HRG3-���4a�F��R�)�́Ld�%D�px��UҲ��g���6�]�v���X_��TT��� o̘��tj��N>6��,������Ҭ;Ɇր��;C�NI�JQC�MOLB%/߽���1S�X%W��]�t�3!�J^�\k�c�Tum*���N�O��d���� %�C6뵅�Y��$�q,�d�9aV2��K7n޺r�P܅#'ܪ��z�m'K���13���K3�[�Á��۫V�n`8���O�c�4.�J}m3j�����q*�p���g�v�޻|%�"����s촵�}���-��ꄢ���ny|���ۢ��S1�	si>Q��0V�%0*�(�+���g�\;(c����9�M�8�q �"L�X�A�__^�[y��8ux����.\��/�M�1�E�Z�P���,U0k���D"Q����8��,��#���{���8���܌�<H5ܪ��`cg�kwo�DE�8#���Y�E~����-�6�D�g��3bF	�!v���[*W�yz�6�A�b;��ya�4����s9d*/���W������Ǭ>x�����R��| �R|X��;w�I�w��e֋/��"�#���}�{���4.Yĭ��⻷n݂(��_�%H�Β):��A �pD���3g��w��]p�CX02��7��V
M	��m�\��%הF�g�6��޽{����s~.�g��a��q?APz��Ɇ8cQ���!��q2OF�$K��Iuۂ������aQa�7�6;��].��
�^��3�a%[�2���Ob�o�j":%����N���&������G���W�������O��O����/}��'O��j��s@QRy����	ߙI�����a@�����Mm�{�V����}��:��[���?����k��+�~u{k��!-��k|9��NTu	XU�����p-Ԝ�"d[���I�89_Remm�m�"w_�C�Xx��ޣH� �S��G~�B��xH%���x:vCp0V9h���˥8=��I��+:,a��~�,���N:|��i��:8�~jj
*�����O,\�|��t��n�m�K`�z�k<öc1�(����@M3&G�7���<��!R��K��tLK�9ڿR�~T��8��ܹ�9�Jp]W��$xO*u|bl�Q�����'N�P�i��(���R	Y�8��s�"��
D*�����|`��H�����l���Hi�W���+>��������ţ��6�~gP�ُ������O��kD��C��� ��(�p?r�(��]&�& MF�]d�e���_������������ӿ�T#э(�4�R.�T\�*)LM�B�_�+�^
�A���z���[U���t�;oׯ��H K��f������q�8��Xu�j��T�.�"VU3�=`?GT��*�`����v�a�L#0�c������봮-_�k�p��S���4L;Ȕ����]�L��h��+��A��?ŶR�
,�婪Gq�l��A�MIESj� +��@Mjc�~+t[�õJmBMagt�Z�19C�m��9�>�Jh@q�X�K(0#"��H����\���	��JG�^� {Cਸ�:v�3yksݴ��ego��Z�c��V����XMɽ �<�J����v�]}LE�L2IY\�cc���R�^x���eE':N�3��maR��L�����[^wm��.�%����������#�0����$5؄��D'��b7��K]�l% � u5��(�uP���e�0Ͻ8�)�ZSռӵ����;�:��,:{��n�jzy=Qӝ��0���]�-`@΀��t�TvA�R�kД������ӔȖ�f��q�b�
t�0�iu��0��C�[�ٸ7���~�E�����fa�5l�!��$p96c��[ `��J�)�� Ir��%�&�	�4�~w�ܹ��ܩٺ��[���4�dg�����V;˴zy��X�����7N(�Bl3��I�9�D%����G�|�3����N�������F�ݠ�K��s09@̙�Y�Ț���\V�0����Q�C~S3,���T����hf�I�Xo��v����U�
��o������|��Qj�e_�����?�'{�.ߑJxE�
�Ν;o���W��N	�bw��V�lo�C�3�eֿJ�ú��V�S�J�8u�x�a�(bx�r�!�ҔG�#��0[1��,E��Rlquo0���c�kԦ3�b�o�9.�R��u=���̨����#MF�@���g�J)P�X�*��=�Q��p(ݑ|q6��������LB���,p1Fb�G��b8�?aN�^%a���Sӳ��zE�������<������ݽ��*e��,M���#�*��X8A�8��~�ɯ�ݿ�O���KyD��[�X�REQ��vo�a���_�;��ɓO����/_^^�YYo߸~��阿�[v��V+Q�Bݼ�`������d�fQ��~��Y�������?~�_��׮^�73�k֯ݨn����ז����Ca�B����OY�/�����������^���d��JՒe�i�����b�db9�)u.���ُ-�¯��4fcb�G7��a�F�\�̈Hp�P�T��@���`��8�8�睷�:�[3Fʋ��?�8���,�?e���X�*hQ�=:��*F}e_���h4 0�0б떖���:uJ�f):�%oof�
�1�/qF��K�v7׆Q�k�|s��c�O?�wnߛ��^��!�F$��U�LA1�a�h؊��9n`�ǞY]Y2�tgc��Ͷb����(!b,�!A�191E9ZF������vkk�ף�����9>I�����Mb�����@$g��>���?�S�֙����ήihGO����/��~p���>3,���m��0ݡߨ6��g�6o��V��i:U�,S�G���N��Ǖ��}����H�A_�c� �r��o�p�p����>�[�����D��0B�\;~���O<�:�n�J�̲����[��
�Nr)S����-9�<Œ�	nj��*���a�Q��9{z����@à����Z�7GYa�~��]%r$��b?��c���ג*Vs-�7�7�(���f� $�Fآ�~�L$si�z�}2
e	,5��N	�u�n��6=;SmN����ފ�Rk��0����;�J��F��T�O?̂(6�W�H�_FP3X%���LOJd��D3������^�I3�){q��U+�43��a'�-�"i���J�H��������"��4"g�|�E"r)�s�t��~��$�Ugw�����S�cY�<�Ynچ>��~�>>������Ԕa;qJij���`||lj�H�ݻ{w��N�P�(o�#��%�3	�F�,����6
�q�W�?t����$�7W�bU�����Q�G�N��5I�L�����w�AUT?Q�c��(���&��ќg����\���l�������,k4aɬ�njVɅ�mC�U{� ��@l�
�M ��6����}��Ķ>%2E����qV����15ǎ���n�K��I�[�Kc�1菄����qR/�Z�3�����L��dI
ag�ؤ��e�g�&�X)���kGy��,�i�Ǩ�V����ޖ)�Y�?��Dv�^��-?�V�:��֨׮F��6q7�p���4�Vʋ���@ww}}��;��DF{h~��Gw1���e�xN���u�6�Wt�6�ߋ�=��^8~�8ל�����'N�x���|�� :D�K�?������������o�};7R��� ��(R%*x,���]��fj�?vvf��v��;U�US��k�q��Z���D�
&Ŝ "u�����������H��V�a�u����o�/��9�9�y^y|$�0�S>��s.@�@����(�i�N���Jհ5�I��p9���W{�m�O%;�Ğ}�g�s<���:,����OMM�� h�s�8 '�����?�.���C�|��(�{��3�5ξ!a�VN㒭�'�A8m*d�צ��DuHIeN$R��dv�21=�F�1�$�C�|��af�G d�5�Z����'k��{O���mu;`4`{�[kT�'P�P�J�>��p��}�v����jn��� +���fs
������0��v��N�)�K�S�=�hCXk��y�H�8�7EW�8�,�
YU�~�-E
��X��\.�Ax���ӗ/|<<�7vmn��ۗ��}��v�^��N`����J�q|�݆�8�"��g.�Ϛ�x��FFF��:X�:�8S{��l7ӍE)m�I&�%�B�=,��a�{^4�E��V ��Ù7?�љ ��n�ؕ/�ՍV���.|NJ`v����s�p��u�e�qߣ[ �$�EY体��A��e�78%OK�-�W��������<npE�6o.rq�E	��slko�����ޢ���k���������_�����յ*<���a���lm������0Hj���b�X��O�嚎�&N�NQ�m�Hq^��N�mum���}�h�����Wa��UKK�A T������VSiD`S>Ôb�J�dBð7sb|Ǒ��n�rIԣD$��W�IIr 팡*�Nn���a6��a�Q�֖x)k����d�m������l.C�X1D7�l��`��S�����ex6ǂ�\T�����,2��3��'w�э��f��|;�|p� ����u�fsג��\�ȸ904Ɖ��I�3������I�nV��Y���W�\F�iի�z��J�F~],�r��j��k˳�������	���!j��U��0:�OH2bB�����R����m+L�B���7��\� @���3��m7M�Ŝ&����±c>�����w�f2�"��g6S�P�L�5�k���N �6�di���ju�����\>��r�h��v;��j�ݩIfk/���q�n��	,�{���!bb!n��Q1�D�3��v�A`��	��F�@���<�� ;����^��NKAQ1�O<˳]��8�$�3`�|ִ;�@�J�RpuU��d�zsu�^|���K�n�8a-�s��.p�R�(�0X��YYY�o��D�$Q��s����pZ
;	)c0�.b%5�:X��1�f@M`]�~v ���$�L6o��,!��8l&��:<1�%M5!���n@�4��J�R�iK2��`a��/d�圤@���`�H�JC��5���E�a��o3;;k
�\_ы��L�N��G
ֹ)F���y"�!|΢7��J/`��(X��u�ܰ-o�V�_���m`��K�յ��a��)�J��9]��9Q��j��$9��b��V.G���>$c��ŲY���՞.�M��uƃ���&�RQ���,� h��$��V��g?���|�#4W�T>7gT6+$|�_����yx⤯
ޭZ�.,,@�p�����1]���$�M{�S�dk?l�������
�zz�b�z}jj
�CXxEŮ��`��Ѱ^�VLOO���Kw�}�U�tX�(����ǅ�n�������-+�ʸ�OSYj�":A��5<�#Y^6���f+8����4sK�JFT#�Ul2J���=�؋�>>�ُ|�4)G�������ə4���=pI}����3-W,�j��(Աr��O�N�)����*+k`�G�F`�Q$rb>�����5h4���s���v�
����b���x�Pn��
�@.z�����6�U����*-Y5T]�_v�6��t�u-0D0H�p�;v��[V�6.O_�U���r�����*J��\J�}��Z=����ڭ�J��f�p�2��9H�l� h1�,\$���pH ��Nfe�U���l.����Z�z�Z,q�O�,{E,f�
Ǟ9�������$8��G�֮�� F���D0O�لŃ��qf�����Y�M�+.dSӢ�$���ő]�'_�p��B_1W�֪�LV�Z]�:�C����EVT�u�i�k�F�x����5��ž�0 (��%`����@�.��>~�8��ɓX�W���B����m�ʦl�ЉR�00�#�vp�<������Qސ17�%;J.�$3�AX��Sj�CY
�Ձ/�x��&�S�M�9.��d3�b���K�rkp�T�![	�#�{�ܟ��ݟB���� 5�bK���V�ёr�O<�����?�7:�޹crhh$cb�*pQ�����3:,{ׅ�.�5*� ����|H��o[mxo<�$!����'���U�XR�� b~����N�R���DZ�\�ir�da�w���R~H�[�y�O�<���	��>��%R��O��@H+��Lª	���h�#�bx�ܽ{vMLlW̲���®��
%�����+K��ձ���n#/6�3�粐1��1j�=���%��;q�lk�$�p�n��f�m�+f��Q,�T)�kb�^�����X���^���ghzc,.`[D�H<��H�x�)�N@]!k9L 3 ��y���0*r�	���]�el��7��9#w�]�_~������qBض�>�񃣁]�5�W�]�"���%Q{B��adu� ���N����+�''&�f ���Xģ���=��SO�����9A�ll4D�υ��czJ��:�
�
,Zʼ�P+N��0|�7�ä�����ܕ1��yi�y�.�]]�v����V�dr��>V=�� �ڎ����*<�%��2c2�u$G�nA9` ��\n~~��t��N�0F�v���P5�0Q���:��+]����󡏽���iB�$ �1�zQ �8R��|^��<<zdt�<�h�( �
kl���{����]�vu�յP��##C��nw�q��A�'���� r�P��$����DY���IG�Fٲl>׵|`"�צ��M�ͩKN[�)p$���p���!���pj�B�ѬA�t�wNMM�XCۛ��{3տ���d/
,��Cxi�A�K�I
Ѷ�*UQ�Uyc� �ͷ�oE��:C�A|��}����m�݆]�d�V���|�
B�n V�J���m{��Y[��O0���(�.#�����(ӪN�Fn�K�
GI�3�����^KgSg�)I���&u< Z�ii�>O\ p��r��_6$H=N�=v�խ����>w��=h�+�Jg/�r��OS}OΣ�F0��zሺn�
�
��0�`;2Yӱm��]p���ݚ��"��h�*u��ڎ56V���+�c
 i$ �f��h��ɒbg�O}G�2���[� {��<�@pl[`��̑��m�s\�lT*��z��8�$��BJ6x��aX'���o�ybZ@k��z��>� �s�"6�+�Zn��
��P��fgg��*�������
�Ϭ�!�C�h�3"�C#�ds�i"��uɢ�)�mwg�^L�&X���5�0@3�T$z+� [i�.�_s�N�q-8�w��Cf���=�,U$h��+d���o��V�-<@A '������G�rn��b��&<�4UϺ����C/��JM��ѱAQ�s���b�r�Ԃ����B�A^Ht�l�=*�80��.�>�{���fT�+XI(^����;22F���n�;�^�Qe�5�GB�=io0��<���pg���m�Pjiy�Խ�޻m�6�m���g;��iU�刈��0|(0��؏K����/���L Rx�|���p��'�P�g���ÃC�npIt�V��@胖��h�^�V��9���)�����W^x�I3�XX��K�t'2ϩlr �ޢ�gr�(qM�#
��w�Q,�q�VI5T��-�ڄX�X�}sJ��z�:^U�"X{`�+�����A�Ѓ�.�r��F�^Y	�����#��l,�g^>+X-5yd��[mK�+����Y/�����E��+�m������NǙ�<�o*�/h��X�d�9�ds�n��{�^>��k��֪��a&
��۩��)>PQ�q40��].B����&rY29�X]\�ػ}����`'^t�X��DC��d�ض�	��x��OWV[R�P��$^=��@����Q��!�3YC56>Jp KхJc.��0`u�jeud|���m徼��x�ײ�w�*8�of q.^���t��^�30�)����FY��5�X���څ�'�
}�G��`�R�6[`��E�;��ȡ�y3���6�_*�U������c� ���׾�:{��+)�l2�P����1�m-�V2d)�f�[A�u�F�kw|�����;��S��W�\_i�StN��Y[?��o�����[���|�vli���k����(H3,�(�P+B~�JcM�r{v�ھ}��7�}�������VW(8�o�Α'���Y�ˣ��|\��^d�7	������f9H��$5L,���.iv�S�T�9�C���@F��=�k�-�ny�ӧO��j�
ESS!����0Ōc�&�2����O�/�b�c�>�c� "mlT����z�u���z:/AaM/�����n�kۼ�ɖc�1�x��}��Ul��%�I�2j#dEX��e���<�uV��o���n�o��	A>Qڤ��C��n��M;�)A����｛���"!����fl�)%)PA�����&E!���W��99yev�֩�5sY�զ$:�G�����fko H)c2!��"*�t���2$ˍ�>I���c���qG��)�!��t�Ce%��H ��mR��4���V�-������:�Z��z���`�se3Y�p�4 �-�S��T,ra�c�>���d2�&�;�T�p�N"3C76j�O�y�����^�O���V{h��):Ĉ`��}���~�����t�I"ow�]���Agu3B��>D��#c�C#��2�ϟ�,�b��CG��~uqq�o����_[��hk(��� �<LMM����:u��C'���:�H|��A�����}5�|�[����Ͻ��� 0����,v��;8���.E4�=�M��UՄ��e��	� 03�b_��YXX��§��2����&�o $L]�l�P�
r� $@ۿ���{�#�����rN�)�(8z�Z!�|B�t�}+�Jp��fszz���$<�O�K��JY��!�_��=�$;~�j�s�sT�p��n��С�o�9_oT�����GZ�)�8�Noiu�Ym7jMX�`_�����Ӟ�:�Rձ�,)!8��\g�32��\�T�t,��+kSS���I��%^�2S�U`������$t�����,�XY��AX�[RD�_���Ǐ���]"��]Ҙ��Z�'�#�)�v��p2p�'�N}y�zu~��a���ڕ��nu�����˃HԨ�VdI.���y�XO#DKF��{���X���~��Ô��ui���}˷[��5CTs�]k�jhQ�+0B�(d��!�tIT��7�*���-_�]Zٸŏe)6��ӕf��2�N��C)ͳɘMJ8^�`�{q�&��z��{K��J����~Yq�/�֫k+M�<�s��<��Og��/_�{�i���qF�9��q�`n/��_�@�$�7���=1<~��^EN��+���Xk$~�)�׊��\ھ�#+q|���`I��H��{㮗��%$�&��E.	�-.�A
�ng}�����f�L����!�AceQ��V�ϖ���N=����Z|��'�vS�߆���Q�(���l<
5 L�v
`ѕl�ت[3.����~]�gN�ʂ������������=G>�+���Y���gϞcAT��]?��9�
Jgr�".J� 65�8�O�%23����E#��؞�(��}{��~+x���3`���B,^�rM6rw~衻�y�d�_��?��VK�~3�'� n��
�-�
�y�&�@=�	��{(cL_����u��������@	'������Xl�:rf0	����~�K�B��'�XX�
�%�Q���I����,�	�g��W��u��	`o�?�OP�U8ޟ��v�Э�l 
�6��V6�� �F� 0�w�ry��޷���$puY��CL8 ���R����+!���^����e�y!t<�k��n=v|���A��+���M�;�z��8r�g>�ȶ������$n��q35zt(8fj@0T�5:��"Rdm��2��ʾx�PV(_��E��0�a#�w�V\�%I"f��YdC�Ú!y�갂m��
w� ��_赕�A1a�ܦ�K�K1@TD|��A �e���ݴU�e+.�RK)��ǵ�k�� ��ɴdD��!@=Uv�4���K�aʬG�
K��!��*������x�jɏ�`nrF(�������i�æ �tt�bb��'�Te���	Ls����8�m�*�%
����B��8��"�5���/:4u��tk�����޽�4�#���I���D�בƳ��������b}�j�*����6ٜ֫��g�+�kq\��	�߶c|�X��ع}������ƆG�GG��G'FU�\z�L&� ��������A��)�7�ߊR��+��>��c���z���V�^�,���7��8,
��jL�{������]#.΁<xp۶mo��C�B��J�)vj+��(���o@l���HBs�=�I�A:w��������5kf��!jJ�c�v��()���r�U�-�;P��612^�VVZ��Țv�{�i�M�LP-���	����"n�n6U�
��9��u����HJ?ˆX^�N���&ǘfR
鴝o��X��L!1��
�$�'�� Mr��6pUc�W�K+�/���|9�7�s���F�	�^]^��o��r�Gw[ղ�r�ԿsϾ�}�2�J���3��)zQC���E�npC � YE�����Ç�$қo����f�;�c���W&-��W,:m��9��p����766�����O��ѣ�ՆRb�S�l-��Rg ���G�&'��V6b�{if�q��5��Z���A�D�����'&v�MlCA!��˳,#�&�C��������Og�n~���Q���q�G<d �Waz"�n�q;�����C�12zĳ� ,�Df��q�+�JeE1��vk�sg_��a!J�.�.��&2�rV� �C'IG���Wg�D���|�Րy�������ʥ��������|��Ս �۾���m�������T���Q'Br+IS��G^����XA��19�GQ�I�������kw;žܘ��u��L�������z�۪4��F��w�qG��㞥�//�\�QI�qm�ݰ/���*6�;[��-P8�k�
o���޷s�?�{�5o#v6*����N�qbU��;�:q�mw����z�{O}��0�fs���a�)z�kKai��`#���c;�#�d��U%�;�w��J�=���铁�8�h�4���٫����������.#�B腰�����m1RԛF�@��$$O�z�iTt�k �ȅ�:�����X�T^~��ZU�r	�*���Z�5���L�_����/��|���:m�� �������AHd)߽�t	o|��''��6l4s����#�VVW�Eɼ��1}uq�R)�'�(�6:���|��?Sow���-��9.�l�	! U���^����,���X���ݡ���;Fc�;����h� eu�B����(l��ѡ�ǎ|�㟪Tj�.�؝�(Ē�[n ��I��m(��� ��B�P�xȉ g���r!��뮻$E=����++�f�Y�t�nwl�}�ͷz��S�0~������46\R�l�I�&�ޖ�u}ºG"�,�
������_�xq���[Mîw�l�ᛜS�"������8a�Z�T٬3����.�:���}(L�H5�큦��&��)QM}��X,NNN^�tiqq�V��R��(�H����u"�{o t���}8]Kq� G�p��v�\.�o&_xW.�b������X2��_��*};���!O�Qi�\:�C���1&@,1�PX3�,�=2�o�=q��/��/�ӧ��c�=633��JʹGc	�A�c���v0<�cSc� ��k�7�M^���?84���L	��)�B��o�?�"KgO�OB>b�1����m�p%�<4��� EL݀�������J��=|�?;08�
��f�V˵|�W�ڴ��;�=���@?N���!�1��W�k6'O��ru��ޝ��S���w^�|��^~���w��v/��N�Eb"~�1��۷6�gϞ�;���;1뫍Cweu�̹7vMI咊K<���˄ֱ�=��-���ԫ�����F>�Į��Y�4���͍�o6q>��)DbAS%n�AS.b�5��]�m�ZY-����**(:|�!`W��9-6�s$�7��MB���	�7�B�EAb(Hx�mZO�%iQ�%���J� ����z�:�S�C�����[��z@B����|��EZE�.|�F/_����|���n��b��d�� �,���:�.�����}�c�l�nn��\6�gZ�9��s�\���nh���J/�8W��wR�e�Ν��.sqq�
G��Ҫ�A0�T<n�6��ێ����#<�k׮i�T��S$�g�4����I�JF����D����\*�>���kw�3iv�+("�`���>��eu*���k׮]+�|7 ���gW�R2��h�K�?Q ���@b!1�B�b/��\�`��P���������ox�v �P�e��(��{}�ȋ%����f��S[�������x
�"�a��'���y�$���"JS�W ��X\&�2��n�]�։C��������+KK1���D��o�\�/���n=v���ν�p<;�A��q����V�x3�8Z�>��O��WԽ��0�:�4�h��%�sg,_0��b�f��}滿������<�t,�򘥩EVUc4�X�b�x�c��$�q(�QluQ+�_�w�ٽc��m���������+�q��W~Xـs���/����;�}���/\�,��{�	ȇ%H߇���\���a9�2��	��m�c˃}ǏU啗_����v���9y��ѱR_��j�o�����_m�99�o�΅���k� �� �z�Ei�0
-���J����.�z�N�4P,�Wk+I���g�����^}���Ȩ�&#C��������'���g���o��Íz������� f������Q�3%U[
�c���9ߍ�h��XN��?<:��O,�����\Y���';6�DQ|�г�J���O�џ�އ?����4�z�T�C����M^�%��M�ф\���q��}��,�~򵳗�._�����!Ҋ��	�F�j��_����Ϳ�Wy��v�٬!KG�1/� -�l8����&]?�s����V�՘��ڱc�W����o�V%f*��5U���'�}�7����;��qb����+K"V����Dq��Zw�KPD�e���eL���U+j���Q�m�K���7�Z7�-�|k\���+4dE\t��-�m���h��'�v���}��߷���MbRO�#	&P�<�1�\� �g_(�H�����t$5��lw,Z�['�a1���Q/"����Q�ɏWcq-/��>���s�G�+�ݤ|�O�w !�<y��x��05������0=��Q�{ˡ��P:���[�k�'HA����/B�g3y���<k�F������s?�s���!� �	q<�fC�q�w`a$T4���4*E�uD�KIhT���P5Ʊ�ݹ{RPd?�%F-�=fs�� H����T:N�.盏=��O.-/��4�m��D5�F���#��
�_)�];G3rXԎPv;J .TL�����;���<����A�{�~�^z�E�R\����2�г��K/�0�˕K}�Ã�����n���j�kK\,K���:V�UAؤP��~��;v쀸P�11�a�R�ݮ��3m�=2$DLq�M
�\"�@+˰�L*�F���0�Z}}yy#���f���c���؏�{*OB�=�#�]�"f�deimr��Cާ"gy��F�'�x�qJɸi\�TA�_���c�x�-Z��"�Jm�RHE���(l��a40B&��[DuE�"j���z�=����&qr���,�j17T�"���U�+�3�(�x6-����������Q�X\�L��h�^�RAX�ŕ,�:��s�حGo?()��
�`��A(�낳�l?�'��5���.��_�\�b#�:������Ú���Wi"(����h����4}w���{��ۏ�m#_��w�Y��UQ���#�NI
84�e��=I����ǎ�V��O�z�R��a²�QF����8m�J6d��n���mTj�9�&�y~ҭqT+��	�}�r{<����ؓ�P�a,�`�����G���ۮ
\ǋTA��+$��׆�Q��s��ټ�����G?�ɓ/�Zݰ�(!�9].x���u��&8�c���Y�'`�%+�S�b)K|}vvi���앫ss��Í�E<*I`�����O��_����������T+-��G�{�S�X��WŃ%��R�B���oA4]�Z�}������P�\#��^g��z���R�q�n����/���-��<<���=��V"4k�F��Q�]�	�K�5��T�(F��&X[M��J��ӯ,ֺ'/��.�WM��)�j�s�4:�re����;vO��g�wp���o�B�.k㛞��:���Qrr��Gp� u�U�$^שw\/������?��:]�uNNT��u��+k* "��v�_����������烷[��(:�� ��U$1c��NY�?�0���MOp�ݰ���x����@)���c������&�Q_V��'��H_���CZ&�ꙋ�Gq������<}�\�}-̱��0^�)��C�b�v?B�)`�0�<4��$ݠ8(��Is�_��O������奪�+&6�q�ڹ���=�����O�������׭�ގ�����:m��xZ|�G��F��݉#��+9`�����`�9��铯�unvqa���5�jGH:�v���0�����~�����Gﻯ�ެVΞz3�-Y�4:�k?�̡fw���b�vC��*l�v��2�ԁAt/����ϝz�]��H(�)�(��.V+��k/�������X/|�m7AT���z��-�>���.�!�7�� ѻ���Q�+R�x�b��`�l_XX������L��L�"��<�C)i���- ��F�I������я~��>,?E���͂��� 
:����5�N��v힂��if��Fu}a��p����8�+�;�ب��ME� z��#����#y�Hx��5Q���~pG��6�l֠D�O#Q�SJ�g>22B9Q@D��Gz席��[����z?��=��5}tt�ܹsK��� �Ʃ�)����(�����o7��ۢ򮵵T/� t
��a`�--�Xl�^8v�n�q���>���Ǐ�r��:!k�����{���b�/�ˇ8�<�\---�^��ȋ!f�!
Fm����w�7�S�6�B�P�n��8������r�͞mج�������N7�8�(&�xN�ҥK�����d2Y���Ե�b�,���*�V{ht�9�,(�u���*�\)g�SM�vKp����aSTF�jw���?��zu��kz�趑�8 <�q���7:T�ԯ}���z�d����k	'	�3�E����v���m���Ɯ�ߟ�;p��e0#�C��".��Gr�4���{Ҍ�"���Ғq�I�?�N	7V��T72:��4�|s	b���­��!@7����u@��a5B�FbN�qX[�D��"튫q	�-��������>|�;�0��QX�-1�ĽA�*� )
�2���߶�T��ǿ5?��cw
E�
d�?�v��@A���ٌX	� $ \���I* .�P7���[���\��������] 	�#++�6�ةi��E��D�! ���ⶂE���W���Q����SA��ѷC���}fT	E��Y�<����TdS8xRp���&��G9p�#׮]�z�*����zQ!�^�Sm�Ķݻ��ݻwrr����M�]Q�l'�9�d%��dY�V:��!�&u�:a��$��a
��tj����G�T��J�S�ru��j �3~��?ڊ<{Llr���V�DD�7\���%S�O���w9��=�G�\��a Q�ip��氜
�mw\��E�DJ�O�'./�)!|���s���=��r	쵑���I[���]��Hu�����A�'h)�0���O���h�riimM�]#�.�s�~��N���^[\^��(�p\Č  ,�D��<�vL0��f:����BN�;9����/�}�U�Ņjݵ�Ѣ+f���I��1[��r�ɧ/^XX_90!er��R%`\���U5� �D�{Fȃi;� � �$�(�f�Ԍ�^\����ʓ/����q�f�AFۍ�V+E����*�+��:����{p��� �$��Ş?�g�}�0 w��0=-dJ��\j�7ο����[Y�ZVQ�f��Cpku����b������J���
���z�f7t'�zXܽ��
�U�4��Jfd8�e|��;�_��}lu�Ip�l��# z��l_Y�]�8{���{n�;<<�m���y$8fL�J�F����D�i���@�Q.��h����g��W��m�!��b��tU�'vMd���g_|��~��>s��[�]:�j�_C��2�q��C�d��)�mǋ���J�gCxt���J����ZǲT��B�f�40��^��c�w��];�������I{x2,�'�C��~�x�Ú�da�'1�\��oO���������eM��`��H"F�bV�c��6�I�f�>���7�>|��'O}oyyy�<�o�B�������Wlΰ�0�+�l�\i�ɡ�~��QW��:<��i�����L�ۓb!n�B(IC��@1�N�Ѩa�n�hF��pr��������UP�Q��ڵＪf����J�R�L*�)�.o&��5�E�M�F�pB+�į��,�[o�����4u�m����0�׎�g������$Y6�R�DL��n�C�q22l@�Z�z�E8!}�7���+��&ѩ���w�3�8{��A.fƐ4X`�<�裓���8���2gѭ&Lu��w9rBj���\��g�y����d�P���iZ=�~h��<�� ��Ω�n��tP�̃{��e�3� ��.2����ҬE�$�Pss�MbWU�h�\�O��p��ZeMU$X��|��+�����PB�����z�< Q�c{���8%N�P65V�
I,��LM/���v� �����%Uu}����b.�rl���lĂ�={�lJAN�m�̔F�>�a�kK2�F�Re*Q�C�L�[�eqey�u}����h�����zׂ�&Pu>�b��cf�C�tCH��zoX�s(�g�H���a��dr+k������]��@"�8�󲤿s�R�͟
}�l+��Lp� )0�䇲��OĪOo��X�oJ M����V�������7-ɢ",�m򆳩qQ`C\@h�K|��HB���	���ą�$���]���Oĉ�O��!�)�'�j
�˄�"�l�G��{�=z�(��Á�S�)�F"x�r�ڊ䴰%���N�'1%��a;#��Tۇs��VU�X�2JRO]	�����u�ty�E��,6`Ho�;&I�ôT�ݨ!�vC`��'\�)���KˤX@��Xl����a��u�D�P<����:��^�%����,��v"*f(�����?0;י�|ɏ
W��6D*����k�|	� ��&��[N�Ƽ_o.�d��p��-�A҈9EU��r��+����.����,.��j�E>����At�Q2U�APp���c�%���b�(&XH1�|��dC��]�Ċ .7"�we1)�Ku+۟	�p}}}׀h{v�kC�,| �[���a�4ԋ�>"L��F�4ʰa+����.��x��{ B�NoSP����%�wK�u?	�������`}���02�b��<� C{O�{\yh�4=˦�Ƕ�\y�P�����bԅk�9A��ϭWV֛�֐!D&�r����!�4��z�#*�����nTױ�<f#5L� �I!��vYWﯮ-��Tm�x%�4��l����ߵf���'ma���'����3��t]�8��D�ARLI����kDE�����Q��J��!U������	�f�k�V2����u�v�>�jN��B��W6v�#s�x>�%K�l������9M���dr�yT,��֗;�3W�q*b]��,��ʃssW-�p;���Z�֯F���5<0a�4(X
��>�vpG�{����*2�����_���e0�����Z���LI�����ڵ�y �T�q��Zm������µ��L�+�\�^n���2Q�B��?8��1+9�z�677W���d,�&ƶ:�t�5=.��NlǮl@�9`6��իg�8_P*�e	3���,ixN��z�:�6�oye���+��c�gΜy��9Ve"ℴ�D%�"b<t���4�N�����һ��^�1-�o�$�Y(����#3%M�|H+!(����!h�n��á\�ͯ�w^�;�����/!�쭢M�T���b����|�}��ly`8�-��<���J�ө���� �8y���˗�M '������h%ÅS�
߼UY�%5P-��g�,..����HQR1�@�N�
�����ԡ�6�2䈱rIt�#��1��F��558O����F �!x��$����7:�F "'�R����f�ju\d���q��-o{��{Q�Qe�5�TI�����/_��{r��m��
^��S$D�5���h�Ԑ`q@@z�����?�ذ�=[��n�n4� ��������5~"���B�'��l
�	�Ƒ�A���<�t�Q�ybtpt���0%:1�Ʌ|_3v����/_�y����?^�9�P�w�h���T��bI�U�M���U�=
[�������ߪE�D��;����j��A�1N�R��r��ӳ��G➸VЀhL����$.T����n���+��� �,��eU��َE����)�Hw�<�7X�$�Cf��*������c%y805 �>�?�w3vo��V{m�I�`��!�C�!8� ��L.�\|o�� Se/8 Bpb��c��*�|�R)���h3%����7U��I���f�ީ*�-���P�k9&�{I��!3�YH��Ѭ_��X��Z���D�|_��3�\X �QBW�v��m�}C�Ԝ�%��*w�u��������BT��k�����)ĝA
����I�< pԮ;П߳w��3g|/o������E����g
}�L�H�6�B�����+���d�",J��}���⤿��mb���/YAW�$E��V��ܘs��eNI$'�r�2X�ܵN�	Q�$��_���Q�E��q��lH�Y4�@�%t�X���ݲ�"�ן�K�9I�t|��13�c{��ꩱ�I|"+��t�>A [�`[>1'��ҷ����<V4 �pR�Ū2�N.b�F`VT}ݪ���"�U�4�f	. ���	^19�|�@x[���uC/r�Cd����@��<Dn����g��[�H���YV-�P�G�e5�(�d*f�lŵ�5)��S���w�������/��j��3�˛Yq�R�{�f�iȞߤ����w� dGGG��GU=/�m7������,�	��W�\ �	��m���8ő�l�~�Zࢴcak����a�����2��M#`��l�m{]����'v�v{�ږU�Uе[�/�_{���U}�:`�=j��c�tr����!ĒW��M�ˁ9nV����z�i�9n�޶2�l�rÖ[	P =�M�A�E��3�8qA�٩5���v�ٴ��+�vo��OxF��J�i��"?�ϝ��/�r+W,��3 �Z�Ɣ�T�{����x����W�1MNN�ڵ{��Ρ�]W�����A��������̼��+K������ �9�5p᝴���7��;Y�Y���峹���+++��O�SF?n ��M��!�+8y8.����J�w�^Z]C�0�	��yQD��¿`R����꫔������*��K)Δ���Tn-1 ����� Q2���W3fr����_B��O=��׿�u�B)�n�F�E�7����;��a
�R9N�R~�
�:!����I�C~�y�g��O}����k���=�b	U�=p�(E�w1`�*,�AP�U���Qeq߁	@Q�i���%�*ȶ	�1g7�k3{χ>t��aO�<��(��f�2{�ʛ��,,-��ʱ�M�e/,.-./�Sصk��@)p�ݦ�wA�07�N+�������;�kvn�o���5+��f�|9���R���aN�i��� �t�x�\����L� ��X���uD��OAQ�*���!�E�N"Jz~�̙��F���v��!�&A�0UJ�:u����A����2pe�i��$x��yr��{����?-���²��>vC|{�a-{���ׄ��xP�*e;�����33}�����oo�^�>�9�pb�٠9���l	,9�ࡡ!�j`X������SE�����:��a�d��?�
c1���Ik�f;���g�B�ã��a�h��.FdHi�e%�h�y�H��ɠьlih���o�?�|�L�47�MJ��{"?�ָ
�7����w���4#D͌�����D�0U3@6���4��l,���s�z��E��������2�C���צggϭ̮5*�������<��-�]�����<j-\:u����D�����8�f�c��$�f�ąl־"fF�t�tE^	|+cHz�rV."�� ���s���#�k�/��W ��uz!��H��͠��Β��*(�ĸ���:a-��s�B24T��K�`���5U���H�F�NE0�������}{3ל�^�[o���'�FFG�6*��q�=�Ŕ+q�`�c� lZ���F2���w����[�n�W���ˉh� b-��V fr�U27*̈́S�R��9!���F@1\D�H�n�3ʔ�,hv��.f.��GF'�M��lV�t;��yR$��esA$��v��-��f�r�eb�WԶ�x!8ဉ#c��Wd1��%�
���}㪪����9���UC"���`���}q��߹c<{�T|/��	Ƣ�[@���!,�����zʱ�l�^���؝8@��b?2�%R��5:u�o"D�by�80�\ԕ%n�ԇ@�Êy<�
�H2�DB�gJmVrX��1���K�ҁN�^�v�V�-M���X���kn?v����Wgf�8��Tݼ����@��w��6�ި�$�~��EQ�X�eef���GM�!D���\\Wq,K�,ɑ�f�q 0� Z6�,2��,�����^��S�c��H%���˄/e�9�ވpZ,�j'�^=��xQ�{���zqx���� ��gg�����_��W\������{Nܧ� �q���;Ҷx�a�}~�کW_600 Og+�H�/:W$��H����mw����"fp�4i��Q�V���A���ڕ+W,�߱k���X�rOt��zG?�۷���Nrzz��q�Q���7��gR�l��*HE`��T��P�<�򉗗������ �i���!Vr6[���C�@p�p9���7 �BH������^�R27B�TJEoҎ8J�a���!"T	K�b��J���A�D�5Y�t{A��K�>}��]��]��� �N6���,�c)�י�^�V뭡���248V(���|��k�ĭ/ר�T[_ѥࡇ?����[;v�aa�I%���z���������ڶ�%U1�4nn.\Y^d'������k�f�ҙ
���`T�%5�|���w��/<���e(�m����.j�0���M���"�GC=>D5H�-���Q�n�ubM�E�h=T�:��]P1�!����P.IDw`������F�� �+kL���/y]V��0uM������d	I���6�b*c��e�5������9�j:��������3�<P̿3j��}�O}⑏|���Ў��ʟ�ٟ=����]{l|<���}�,(`w�ԑc��F�G�+�:�؂�{l7�q�%�`��;2a�rYk~%=���.1�D�-:k��I.RST�,���͈Ѣܓ�f�Z�}�B�t1��ˀ�wqc�)�{�4 ����ƹs�0і��2aC�SO<;�$m��:#Dm{��ޯ���h�ހ�nܼ!���b��ni1q[�8�j0R��w���o�.�V���K9Wnce��������F�,m�ő�C��q�pa�����'?�����_>������w�nKS$i:��h�4�B#G�`hY�(�kk+�������+�,�*J�ĂTi����9�C5��CGv}�c�t�����vx%����ŋ$���l��{�l���E���3�k/\[������?��_�ջ<'' *�L��"��[vcx|�W~�&���s��7�;vU+-ܫ~�
D#[�+� *�ڝ8�c�������!��!żа|-?x�C~����Ŗ����D��D ��P;�=vx�?y���m�;w�u&gp�'pہ��<8*�ϊ&�ACM����}q]�������plr����ӕs��ɨ��mQ .E�3y�n�O��_�R>��ߟ�Z�P_��\�&yoI�<�Jw���D�/���%!�v!��� �8��C�./=�u��|��<$��CnhD����?x�q������xc#1 ���f&cllp$O˴(�(!�K!����ڽg������3a�c�=L��EM�Պ�ş��#;'������]�`� �B��9\Q��K���P�5O�{�W'����߷�'����.�[�\ ��:�����U�0��Vg��m{wm붚ݎ�}�.A2m���f�� �^,y��5��K$�C"
E�Bd0ʟ��gwO�x���4���#u"�up����
�s템�w��T1_�&�Ӎ���Eu�Ԝ r|�(<�@���܈�6�=-
bȔg�a҃OEgH�N���4N�B��+pCQT�>M7B�xP��P.�||�&:HC�e��LN��;33�74�N齴�A���oGF��Z�Vk�S�8r�\؜��c/
��X�~
���{����� ��X�>8�q,��,5�6C7^z��z�>9�{xx��1C�!m���ѩt�i�:%s��su��C�$%	�OQ�7�Ǌ�emRѡ�1�s�<v�����?22?æ�ַ�u��%�j��-�䡉*3�qp�CtU	f���B(�I���`��x]&,���ujƣfN"�v��q0qg���6� �ϑ�������ͭ���,�^;�־���5���n//-�:-�4[_�'�������'�o�S�ˋ�v��c�W-8�#G���8r��Ο��6�����2+KV��3Ԍ���̑x@3��N��
q�V�?	4�0X����29�_��]�Md�"YcJ�aZt�\h%N���F��9l�0�Cʚ�44800 Ɛݖ��h�!��Y��i�&D���7.]����Ͽ4����!"�}QR߉F�;O"Z�ش��9��q�
�GPa�A�F8�0����;��Oy�S��f%�L�q߽w�}�]	g���������=�m[�	������:�!U���Tx8�F��]X���!^�c�d�i1�m��Ǐh3��E�tmsĎal0�TF6KY�;�~"@��&
p2�����9�ٖ�h$ւ�ٷl�]����4`w�������*������ 0\���Os(?���� �w��w.�V�8R�g�d��u�~������8�-�������w�Z�4XbA�i.��,�:P�X��}���+�+L]��W���U[kW#L��b$���t"F-�mQ%|����^�>��P9��S������+(\����M�jۜ������/�≣{g�z���iQ7 ����Ev .�@p���g�/A���酀,�#aL֒X�4��?��S�~�µٿ���Q�z]^�š'��&���w������O>���/�a2�K�*��pb6ϭ"�i>F�� �am�?F�8��с;R$!_�՚k�����?tb�k߶�jF�bQ��j(��j�J��o��/�5�ʋ�_�zi��IEQ�����`������p.���V��Ø���*`w
��l�2\���3�|�3��Lݗ_~��n$�����(_��ĉ�/~��������g��r����^f��A0���d�Hc����i5q!v��҅���'?��O��[y��ץX�!�օ�vpG��Ξ��K��9���O7��� �#��X�C���Ŵ0n����ko���ñ	8��ھw������g?�3�+�W�U̨3a��"�W��g>��_��/���=���c�㊑���6-��XUM1�L:��
�4��q�э�������&���י������[k��B@�bG ЂdY�VK��ܖ۲nɞ�q�D�����vtO�t�=cuki�v�$!B
QPT��z���r��ۜ����^U,3#��T��2�����9�w��(�۷x�=w}�[�;vV��i9}Ԇ�I��P0�?���d�'y�����v˴��5|_rc��`]�)����A�^�}ݡC��s�����G�|zf���
8\?v`%Y��VVV���~��;�v�U_�� F�*��Sg~���Wj�Re0���*,�$��{q�k�,�!�Y,9��_����W�Mp�eђ*Z�R�����Yx
�� 3Fi&L�q��&p��*҇M�%D1,tl��A�Ww�p�`ee-(��&��r� �,��iR��N�HQL�EdJ�����Ȃ�� 	)¤ڸ�́MNN6�5@�O>�xq����S0���/�5��iC�����/�]��8���i��5n�
$i,�b��p^*�.c|�~�PĔT��ʔJ�]�v�����]��k�P?�+�?��{���F���H5�h��~���*��Lw;��T؃ �_��\�wb��-r�?�� ,@ӿ�ms�"��P>��p	�Q�+�+�'EZ���Ty�w�MS��ԧ���7��[�����f���7\p�R��V��
l�X����[�mܸ�t��}�����vMiתv�����_�o��u78yr��JKѧz��ǟ|B�d�qwn��������Oy��4���{Y�O��D�hA`�={w��©��ϜÁp<�w���r�L�%Q`��xe:���>����Բ�N!K�oX�`U|@ZAh6�bnjg�R�T-�Y/��\���۽�R����Z����%c���&g4��>���#&u9$lpa4w��qf���/?r�K_�\hX�L� �A�2�'�-,;1V޴y��3{I,H��c�yQS�֪+�6`6��~@:E�;�px��W*�;������m�h��z1gz�hqZ����fa�g\1�D+�F��I��:�����؅��D+�p�<C�KHR��9J�(��Ϣ�+�gO�l�*�-g%Q "D�1(���g�=:77�� ��C����9dm��ɮ��|�P����md����,���Y�9����|�ʢe{���N3�WܷcB/��=/	�h�3�,JF~lg!�s�ײ��V����[Y`��-7�����/��&9	���t��ݧq�������\k��d�8�7����J�3���W�m�ID�W����y��w�����<���=t�U��d4���H�z��Bg2���s:�l��g%�,�I��{��������"F��/�u3������s��}�u�G>t�m֞y�ў�'ˉ�y8dh/�;&�rF�#;>ŵ,ψ�{��X8W@�j�3�=Jӳ������/}����X!�0�w�s�}�~��칇| �r�Tr�]ـA���$E������[A����X�x�R�Q�h��z��L�X��]�ى��ĩ�^��dN@��7o���[������4��9}�\�j���ټ���3�,<	p�̇NJf2;)fB/| v��:���s��r�o|�}s�sgeN�_�WC,��������?5_8��3�F{��],�E�s|�	.�(i��[`��H�s4�fp��3�F�?yj|l�;�q�����>CƘg�y0�A��;��/�e�`|�?�lo�2�r*�>_�~D�Z��Kt��z��`XUV�ꪑ0���ӻv����w����� l0�Ii����R���{���/ϝ{���m��3m�.�K���T0-�>���ꚾ�Y=s���-���ǟx����[o�����G��_��n��eo �vH�����O��bx��iI��e≣G~q,`�;w��j��H9!���qg�J0x��?�a��N'��C�L
韩q��L]�bgs�s�tP5{�f�}2��\�Ny�q�,x@D<�`hz%�NgddD׍��b�ӒIB`�DK�B�/p�+�DQe��Ñ
�A���yG�� �zJ)Y��ںu����Ν;����?�����ڽ�s��)D�[`��b6�����@�iN@�bcй_"\�DJ:b�LL�R�m[��
=�0
��,0��7�}zi���w�{�����5�@XWSGm�����t��,�`5��ՁC�jY&J t���|
@y���G(�@p�n�Dnff{;mZ8���L��ol[��B�ҧ�>�lt;X]���ϖW��o]}`�'?���{�����4*���M�ou��_��"GdԖ�8s�d�W+�L����}�����܉cK�K�]w�*K.ǒ����nUkU��q<���gA39�B����S��<�Å�-��bn��UMUe�q������)À.$P:��C#���	S�F�$9R,�88v�Gt)�Kg��^���F1V��v�<�ȱw�����klb�U�D�`�N�vCz��V��	�g�$�����M�1���2�d�ܕG���k.�MRR�u�f%�$:� k�8��	N6+I8U�z.oy������"�
U�dv�^��f^[[��L8������>�&V���`���0����{�h���'��(e}�B!8U�9�^�w�A��,ȍ��� �� �d��{��>�P)����ݗ�}�����b!�J��:�/D�9����s�h��E�O�]|@/3Z���΀�5��H�K!�B&���
5c%>a.A�[��l:/ �7K�}_��lpLL�t%bLߤ4�}�!J����:�m�bɵ=�g%�	����Ĳ��c�+��D�ΡD��*�%BE��b4[~cz�	Ϳ�7�N���>��g?�����9�IH�#�X���VC"p2���+�&�e���s�g�g������Q��<����v��9aj��w_{��������/�l.]�ť^����8�U0��D��s��$�����(�4��$����cQ�LMM�]�~����vם����'����PǲfM���w�s3_=��w�|af,�%/j���}'H�	Q�L�y߳4	�9$O�CǨ���BD���(lbj�wV����\��{�:UR�=z���]�P0�\{������o����·��������X�4�Ç ������y�e�Ì,P�-�ȩE �}����eA+��6n�|���'?�{��������G�:~�
DX�LV�����;�}��-�_�)6���j��ױ��b�e��g� +A�����nQ�gCQҶ����o|�a��n��?��Է���#�=������n�j�>���������o��T�S��k�T%����š�L��"�4����M�?&9�E�K�m�G�>Q(?�ǿ761��/cq��`5Ed�9x�_�/�޲y���ԩS� FG&����V���&0Qh����%j�a/)��
�W]+?{�1�����������ӟ>��>~�t<-�{����rۭ��{_|���O�<���F������-��V�Vhc�r,)*0r��\"��c���n�_^Z�0��H7m۶��gNHj��|�j���WΞ��# A��Y��������{vo}��_87V,<p��Μ>�āSL���I�(�vߡ��v=lu3mY�g�/��+����*�ڤq�3����igE:
�.�iZ8e���-��1��Xݽg���v�WTl�������z�&�v�$��0�,�'L�J�L<��32�����680�;@�&�='� K#��H r�!ů	I�O���E��x��I��_�.-.�رL�juŶ��v�شi��[�Ea D��c��������/��¸�t��<qdiaqbj���cK�s�,;�{����\�t���i�J:+�n�t˥/�$$-X��9Х�'8=��(I��m�Q"ϙ�~�<
Ȏ�W���XN�(J<h�X�Nu��a�j$�5�L&�Z �B�%�7���
��_�=K��Ҷ��:��ac	ZX�E*&i�T��	t	���.��A� %`�?9^j7k���'��꾽���Μ?�T]]�>}�}��{b�ڲ��)Z_d��u�J~|�o���0�z7�р��b��ϟ�~��.̟߹{�w��6�幅��]\Yn�{@c	� ��#�Ǖ� 
,P�n����a�ZeQ��C�����>Φ�ɞ�Vx#E��EQ�K8�^��#���	����yw�����0D���Xy���Ixf�3 )���m����x�Ȇbv��k]�����YgJ��%�.���%`ap�|��'��6,�� ���X��ugD_9��zSCqJ�.=�,mH���0��vZI�h��e#�X���Qƣ׎X����&k�k���11QYY^>w~���'ϝ9:�^� �P�Б%�p���еl��E>���j=mΥf�2����]���_#S���f�ߟ���ݾ�Ѯڷ?]��J�#�!^VY�l&lyV��rA��a.M�0�'m҃�b�R�K���2o(��� �P��yU�z8v����T��	���/a� '��*L�S�"�x3�	�w]#�9	 #,�L�f��y�xq�di�(D�v�ҶH�΁���JK����5����Fرz1�۰s��l��_�p�%���P0��$NȂ�x�A�e�WUQ�$UZXZ��W�v�գ�n<���M�N ��؆
'E��t�dcuސ3j�>��y}'�^Ŕ\r��C ��#��J����!�oq�����9��?�|����8�я��B��gs2 (&����6��z�0�DVf]@�a�pV +­�LND����ޚ�ʞѭȰ�X9�)�{��ǟ�ܰ��o=�ַ�8qz�ѐm���GJ���=7}^UUX�j����a��q�*v`��3�( ���P�H<'���aFF*�O�����Ye�D�w�u��o��a���j6+uj��=��ř���Lu�αIJ2��8ҏam.�h��;� Y�@O1]�WIY�[>.ۼq�~��o�����f�$����K��{���Ǫs��b��h+�9Νi�}�%���fv �'օFBL�a����衇���Ӎoݽ����W��l�p��-�b9r���?�3�*�S���W
��"kar�\�wcQ����<�n��%�0�;t����࡫�����w��7=;������M
��`uq���)�2u�>���"�J�R�����A�h8��x�1�c^^ԫ���������n Oyfzz�V��
�k�y��{�K�̉���^�5�/�L!��Ce{~\��G��9��h�8��R��;,�ƒB����֋V�v}�q��5#tYCp*�Z]"��8=�|�0>>�oo��_9���w݃MYpp%9�����(��PI�*��ھ�F��hw*c���q���ǁ����礡=L�XR�7X� ��t0 �r�W�yYX�����R��i�u$�_ᯃp0���f��+Q@F_Iq9$��X�o,.щ"��v��q�*���AO�:])#z��!�O���KDKͧ�	 5�|Z{�Px�0�Jr_V ������h��<+J���#:�jЯ�v�|�8q�l޲�LF�?�&~ڎ+�9�d��`���P�ʐ
' B�>?~VB�e���i��P���5��U��K sp ��vY������˙It}q�l��V��z7?�{�݇wm�K�W�(������m�le�����/v�Y�������ū�S��h�B����mBniAi���R�����G�"`@=p]8�bH��fG���� &	b�Qp8����Sm� 
�8�8IֹT*X��q-x�٬�t8ىg�^�Ё���˱󺔕d�Xlc�d�]k{n��}��R$ًl|�K��FD��ȴ�n06�RA �p�����D�,I�+	�u
������+��GXl���l�g�j�&�*U�W$ _� K��q�f��i)2�8���G�8x�����s��mC�C�D
�a��i�*<8���iںc�AZ?��N��;��bE%��I���D(\�a����g��[�E�v9F�f�.N:F� xc��vw�ZǾ��8AT�z�~}KN���H_C� 2��mWcZv�!tG�%��D��^>�����$'��3HQ@��ɯ�~u�A�NB��>C�Q&���Dd����T�`��B���3\[�T�S^�E�� /��@���r9NdaS����-�2��A�����c�<,9Lx�ԅr&�j����WFFFu-Kj� ?+�K��V��4��A�1 ����A�>��Yx�n�<nw&Hl�<Ǩ�P�fʥ\��9��������X0����ڦ��M0��|��6]�Wy+��1�h�6"�Qj|-l*V`y!�L��цBAH�0�%�Y�t{~����҈�a�nx�ƅ��v�e��m~v���|5�� �"�*��BDt���"JD �=IM7pv+��,,8՚�S�,#������
�^���12z���˪A7*Q��1�`�MH�"�
�\/��gH�b���R�ح��8�L]^X�6[�E`���u��p~h�����{������q^��#��?GD��v��4Cꕰj)���`�}��&U�F[������ٱ�?q������۾g�$�˒Ɵ9����ϭ�U3������e`d8,&�PD����:q�y��iJ��	�d��J��W�`�WVV��6n�4:::>���pn��g��J��iU�U�Q��3l��r��*H��ێ�G@$�1B�Ē*��n[@���Z}�������߁[n�n�q��3�1>R�j���p����D9wn�(�F��qjJ�OF�h@#XWIb�T>��z� 9��3j�! �J�b,��;}�C���_kF��d&w�F�Hy�G��%Ȯ� ���(1oe������ӧ� ���.�J]J(pHaF5`��`�x;s���3s����� :4���~�;eDo�s��4�XX�}���i ������
)1�^�:�$ʿ�ؓ�9�rR������RJ�bM��D6�e8ID�aؗ�%Ð9���w O�}R�_eE"-��qD�� �>Eީ�� -����΢u3[ؗdhgΜ�]�gϞ����Ɍ�K�H�@q��ho�:B0���Vt��Hf�\��1{\	�r�[lx14��GGT9g`�ܥ����MfG!%q>���C��g�>XE?��^�W˙�x�]{v_��Ԍ��7��UF'O�0�����}����ۦ�n��D�cr�9�WOy��l,ON��0��U=�QԞ()cc%Xv?`Vk]�i&1�G�H��20M
��MOO�x��$���$
@���]�tZAIx�`�otۘ*�D�|�"J,�r!���;������Ԕe��ILt8�Vl���	��<���{n)Wl�*az |]_9��VWV���/b�0��D���K^�!vA��gb������A6X�+ʂ���a�,�$����G�tE����L���:�B��zݾ� n��� ۷o�|cmm����]��(���,�Jp4�{�`o���/�,G2���LD�I]�1Mh�78.���:5���=�L�R)��e�J-..���7[؊��qL��\.��;�F�=^��Oyzvv����h½gwe�tC��o��0K��@$b>!�h��]�F�h ����E���K�+�T�q�p�P
S���0x��kz�C�o���}�� Rr����P"�Ր��bYՋ`�Aa�l�-���򈬻n#�� @qb�:�e�d=��ITՐExl2/�2��xvt�r��=7^\�]]n�IC�9���X�X3E5#�f��͌��DpZ�t���PNys��O�����DR����$�cOՑrQPe7p�]�PZ��z�N���g��ZM�[��TE��<)X�3!i90�"���qV�$�-"�o�E j�0����`�%��Gs�y�H�'#��s��s��p�<\��o��6��by,����v�\�s"i�1��y������'ͷh#`}�S���+����11���u� �V��z��j� �#���ceUQ�`���,�C��$���i{�Yl�^	�	�[��Lp�]�j`x�1�����WVW����P�ﭔp�����������L�L!�\�HL��z��!d�H��Q>k���[� N��n|��/���Ĥou�Κ�Ď�d�L�P���z`�x�-۵lxn1ia3�B��i*�0Q����U�󥼨a+� K�-��O��Bt�B!W,eqvk���Ύ-{ybp��:܉�/pZ,i��4""0'-#%
!�t�peI�Eݲmk���- ���Ks�V�GC�a�-5��O�P�����-7FUDm~f�g����1��h��E�E�t*E4DۈR���?�!w RaWt{VZ'��K��8�#VtT1���DoVZR�V'�Yv�c�nk����R�)X�Gҕ��#8bV״̩MS��-�M���qNTY�����ײ�,� ח�3y#��h�[:9�n�^�gQڲ	!B2WL�{�n8ez���K�7���_�~�����.;&�X�>���������lճ��Z�ܰ���*�[� �m۶����va�>y��4��d2�ثTƍ�g0(٬��eXU*�i^����k��/|�_��h]�9<�cǎ���Pep���-�i�{Y��
�QV�w A�'8�W���<�Z�|=�ps��a@��v��+�
�	Z�1xI��~��n�	B,w�qۧ��_dsů~�����Z��1�={w�z���gӖ�`������������ƷϞ�>p`���J`}�iZ�K�|`:t`���-,.TWu0�Ų�xW8�����h�?��/�/����CM�*G�E;ԉ���9n�af��,6đ��8�3�� C
�C<9��v�����>�� ;�ڶ�h4�a�^����Z:%Ӌ�V����V� ��M�y�^��,^�K"<Z�v����zc�1W�D�M	���Vql���n��NJ�>�s|�☋UR!ð����NU��28ZK,'�|�v�>�D`�g�;�hl�ȏ���	=��楓0� ��0�����&��Y�̒���U���V��`Cfk�CIƏ�����)�ɪYj����m{�k���p���(t�R(\U��g�p����V�5�oy���D�}�{�?�ۻv�]n�����ѣG}�aj�ɺ����"B�:]�Tr	CcKQB\.e��cS�DU�Q��8L�yM���ب��j],���̕q�@,V�%����X��a=��}˵�n<tCQ�I��e.��l� ܏�6숑}�������˻޹�.��%�"s�>3d���11Ɍ'��D�N���K;����E��m1޶y-Kh�ڼ 䋆��㡰Z&���,�)+�l�|/$o�Vf�����jk�<���!	<[�|(��h�T&�c���S�\�b��JN�ڡb�j�������d��b�Ѵ�PT�,G0����L�(��[v-�],�T
�V��?^�����02�,f2�d��:]l�Ʃ�|&;�2=���d��(v�Hz�g`\.���e��Z�bd|j�ڒTcL+¡�<pf�u���q�����.X~�%㒱.��I��0�s�:���o6���&7n�����&�]��%}ǌ��N	&w���v�H����e��ɭf�!��~<�h���b,aAT�� ���[�����JՐ��|/2]�|��"��0T3�B����M�N��c�e�����: ��Up�LƁ�+�z����ɵ�	V6oڶ��3U)��3�GX�.+*#�Bet��p���U�P3�Յ����¡Ow�3�S����<��G����VU@r�F�~��������b�T �֨.�-�G�6�Vy��i�Ho�{�n�x�����j�����4RNa"u4{@�y?�����XF�Fp!t8��s�V��+4���笠�6?�뢀�ʡ�$`�^Їg�a�l���ʺ�v��Z3����Z���a]�֬	�����m'�=�\�N����@e��$�+�^�4�_Jr
�53DO���
g�P�Q�gz����X�r��/����_�� x4��V ʤ�\ ����(���<*F���PjL?�������a���t�izG�>v���̐��W����y[����߿o߾V����~�'�\�{ll>�
�?PQ��B��,��v(��c��1�������!i�:�hI⃃'%M��v�}��J���7�L�}�/�3t�-�Vp����y�;ߥiJy$w��nٲ}G�ufMHD&�r�\!���z�����G?Rs���z�ܥ�*`�\V۹mJQ����NpO>����Z{v����GFF g�а��^�T9�&�i�b��ƴ�V!S�TQ������pQ���i�(� ���*�
��˲�{V�k�̶"+�&s�@���j=�nuL��{F��$U��l�ڱkonb��O�|^��ی}��X�|�ȋ�� n/�gv�����R�'0"A�Q�n��Ί�G@�����d���e,_If2YU��0��~����� 2���α5�h	FP/\��"d�p�9}tt$���Òe��4͞ ��Ԁ���H�=B/K���ɃD7�?'���8�D9&��X��H#�wt�.d^a��9���o#I�$�@�T�$�٣^�1fX=�:J/����/�/��%B��{G,������mF ������ 	�^Ɛ%>��V_�L��+�f����8�1�M�,��P2���W�(�ecl|����3�L���6$!���*{��  �#?=rg�8��T4E�5Ɖ%�;9 �1X0����dr3�-/.~�+�ϝ��m���ڦI����p<T�$�9�sl��Wa�a�ڎ��ToV�V��O�	�#�F�����eB�M�`��
�F��������ӧg�	��W���a?��9��k:ܻi�4�`�Z�T����J�x!��/`!S&�9%��>������\��U.-�}����2^9�����Rւ���z�P�T\���Ե+�P.�W��Y�iY�v���<<Kj� Q�u��:����#��G~�$�Fci~~mf�#�гX:
D�xq���R�@s$(�
���^x��Z�����i��&b�"$Uy	:0�������JQ�f�V���B�����b'�gv{@k]��8-��Vk]
��V-'`�ؾ2��������f��2;�Fx�W��ЍQ����X�.g����Z]��I-�)�s�Gs��ӳ˳U"x��0H�(Y)g.���Fű�}����G6n�\Xn8>kY&����!z8�]'vH��q�Y%10�lv��gO�x�����GrL��c����.�A^2�We��.,.���oݺX@�i�?D�
�]/����4/۽.�[����-�ٲ���}�X�>r�٥Z�]��|6��f�R�4$B4�ƓQ�]�q�m��|*�D!�k-�K�N��i�9Ur�͆<�$�J�Uӌl����&eO�UWc�-iZ%p�c"<��hY0TCج�3�v-����[*dq�H�)��:c��{�cO����׫S'�j��v��IPR���*�\��+�d\B�_>k�^��D�K�
s5D��c�o�S��قx٬�}�6�q�08�ؖ�a�
+@?X@���y��۷o����e������	4-Ch�~B�#4��H�=���U׊Ų$�W�-��A
��X�'>�.<���gϞ=~�8�hbb�6n��
���&��}��[�J�{����P1��pf���Vu~�V#� ��I�hR���q���PT:T�j�zږ���_<ݷ]^V|�ݹ}�����ow�p�A�QFϩ��UQenvz�8R~�=��xn����G���:�ٱ��;��B�_=�\�2�|���m��H����L�=�����\�Y,��~�'�p��(*͒�z�� �u2����|�r�$g���Il0E�L
`k��U�� ��c��NᵖT���K@�H�/����Ҭ(`e�j�/�0)~�x�kFl�
��[6XUsf�u���G�����;�nَ�[(�Hb��
-6#�2�l'��"N�q��p�A�+�GA3B�o-���_��UFK��v���_;����H^�Jt
��,����*+�"p��p��!���&4�-�rȼuw����I����-`����r��C\A^4�@��a�
{R
J4�X�� 6R������O�;"3��_{#�2�U.k�ݻ�СC�|kZ<�����h1��kmмL5�2��7�	"/)��fٓ)�����1+Ȫ�P�����-�ccE�ܽ07�`�Vn�u�r��/�|�4
aS� ���ǈ��c1�-����B5@IL~%���xfP����%9a�ޅ�=�ĳL��5�`�A=(Y���3��z6i֎�b�pZY�I�V��_��w�$Xz�����E����v�!4ԅ�c:v����6�*��,�u"��I���p��������ly%�h�aOO��G�~�Q�q����	IDe�p��H*=-�HF�"�l�Ł:(�r
�ɰ ���T��	�ēB ΋��J�����%n�φ��ς��kS$��P��,��d�J��
�\*���Y=�@Y����#�jr@�-�F3@ش�+��[��?���X��K�z!�ka�,:lx�]�!�v� �D��0��>f�`�P8K�ň�%����� �8������_��rF^�jy׋�����-Duo�F��DΨ�j��Y=>��w�NgFq����X��;Q1�K��Pg���1[����o�����ae\O�D��Qh�y��� �A�>��r�WE��|��n���1�ݑ�B9�����mY����� Ƣg��h��ȚfHN0PQcɶ�,�1n!N ���c^������� l��nT�uT�򃕕��믿X�Te7�O]��(v��6�z���@J��Z������ύ�'^xѲ=YⲚ�}ye�tu��2��G�?�Ti����n|�q�25V�t{/��_���hY�����u9dB"���𵵵ٙ�M�ppB$Y�0��J�"�vi-���>�ذ�Q�NWԡ�6�v�S���ucf2�Uԧ��}����i�%�o[!i��4^]�(�p@����1;������:�3�^�6���)Ls��mC"���QC�/�Q�G�wp�Y�����
PhB�"�A��a�l0r��)g �d�zT���O�jl�#���9q�ġCo���e�5/�8��C��v���>���hӎPXߚE#p�����J#��0��Z^^n�Z��F�uM\p�R:b2%]`eP6 �T�@
�G��tf����,|����M۶'^�i7\��ʈ2�c]^9�g���p{qx������dyv�O?��-[6*+ˍ|!����W��̿��м%�,�SE�\$�{�ɓ�7N��f6���W�-l��A����C�Q�~K{���$x�1:E�mw�+:.��j����)t,YE,��}@ۤ�
�4U�?ú�Ũ��P-���gƊ��$C����QBsF�TC���������t��ޏ~v���)Xa�n��V��뮙(��cM�hX��ƲpX�H�U�K6���lTHǙ~x턖K0���u�:~��@�&ZY��1-�gD�l�M�6|�O�y�� �FĘƖ���,��$|������en�67��UQQ�����L���(k!��a���ɑ���4�@�Qq4~���Tݑ�V N��F&C�yԂѩD���)I����W,���)�s��^��"
`� �%d�k���+��	�غ뽑��4#�S��gi��̙L�ދ�a�GrW��z��k�߿��
��buq�g�?��Ϟ��
2N�<l�,$֛�:����Ѓ��S6�a��B�\��
X3I���-DЅKd0�+.�_b�a�s/���W���s�4�1�<�&��۰)��"/%�+ ��4? S��Ȃ�(���L�EX��]"fO�n�]'&5Q�(�A�۱HK=>.���C3uƔ˒�.�)�Y.����n��V���(�� '�1���r�xU�㉲C��r-���`V@�cU�Q{ܷzX�E����!���_a�cbJ�t|6�g#y�n(�%��3��TE�\晴�s��!qi��+�E�s�,�C���Kὣt�ǱC"�OV����������#�A"#�H/A!�*x�u�>횃�I O� |8�`�"��4T��`��G�RP�߁4������{=+���t�@"�nh��8�(l!�~�/1	 _ȳ�$s����0�d�
5(0M�בN� �jìV\��ҡ	��1W�% v,yJ�1�!��OP�m���R��G�%�'��Qd�[KS�"��+v���ϟ�m.ٱ]�<�"�,f�H���j��i����($,�%5��B�O��Ŗ!������ͨ^"�[��
GQ�8�8I�(x��'��=2������<w���=�6l�b��b��s�3��^��7XR$6����x2��|����������|7��J���F�W�#�J��Bt@;�d�,��6<qY�����j���r���j#
a�	�d��X!^���s�L���^�{6�%�i �E)���z��Y�4��~8�\�r!��� �2��|>;7{A�3����KЭxY?�+�z_i�>��X�4�0�t瓱�t����FM0A'{�,�s��$�C�UZ	CG��},�b+�ՂwN�W^*o055�e� �i��e�$����QT4��)��w
����0�B�  �$Q�2c�S}�]X(�Ki���M�v��111m�֭�J��_$�O��"D�ͧٛT�{�N�x�f�6)�rZ�Jo`��j6���7!���P~�h�В��]������xe��[o���!�s^<{\��ܼ$s���О��ȍ��EMm�<p�����7��3w�}�?�AM���C�兏������3�������?�{�C��=�������?p����^6���ث&&+���9�Y�	GA����o�w׮]�ngΜ�����xS�1�f��À%20����
2�Q��,�2"+��'9�0S,�A�<ȃE�Ru�(����
x��\n�\��c���e"P�J3�<�nw^��|������[��m�ǢJ�
�9$��-7�G9�ey�q{��� �A����W�%W����s3�v�ӊ��b��*�dtJD�˱�_�1����I�}�=�^�u'o�Z�3N�U��K�����^�wc��xy�'��jb��jmmy���#����"-���z�DH�"E�c����D��1� 6ɏfJ��ͷ\�g��wwMڋ�W���vLسi�����_�uv���j�1 <�ż9�j G�.�� ��ƙ3�L��ݨ��}���6O��H`5�f�Yb�^ m�G���z�+�
���oZks�N��B6d�g�:�o��m�/�:�	�PHJY�6[��5H��<��gy:�Xb"P)�*`1�$r8�*!�`�B)�C��񜨊행��2 j�K��fKyׇ_v )�\�%2kE�Øն0� +���bҢ
(��
8I@h/��8�y�l��Y��E�B�\��Jg��1eEn�[q��WWሃ��p�������i��,[��b�K������q�^7���.	����.���l�l��,�p��ߪ�a��ض�^L��"���GYa�h
!������#<)xI!�ELÐ�oN��UE����7&�u;}�a���_�� G����>փ�l�H�&d���dk��ad1�,$2^����E`�2�`��H��p��,
87��D*���k���INdUV�AiB�T�,���حHj��6]��±ȨY�Ga	a����X��b� 
El��7�1�$ +�0��0˳Ѽ��6�G�a����Qb8`9����"��1@�YA�D�D��l;E��m�n�4�iB�x��`��(�� �`�8�L��F���"�E6��L�#�D��Z������E�q
9�q��#�"a���~�A=��<K�M��p���2턴C�1>DC���IE&3P��Z�ȕ��Ŵ� �P�������%��qDvmm���eA^]^��x����^�J�r/�x�@���I,X�q�w��D��MӪ�;Z.>q�āh�,)�X�6���͗���c�C��a�O c^|���S:AzЇ�EQ/&M�p`(�PRD.�U�]�^�������c]{��G�弡S����fW6L��/͇��V�!�״��� �x6�;�: ���*LA'�nK=��C�T:|} �G�8a���� ����a����>U�e(���� GFG3Y�����+�=�<!"z�\:�>�be�������`����Gq�3����O��6]v�76J��g��������ad4UՊ�r��)
���~T�ǵ�ۛ�����,py�O���
>��b���3L�
������#��@)%�d�۪��5e۶M�vH<׶hȃ
��|?��S�`J��w�����\�������4 ���U4\����s'�wڽ̲!*�z��m�V����	<j�d���	%�	�C7�m�Z[Z��7���w�}�(H�b��:����͏N�V��lH
����fWU����3gN�;U�v����V��A�4ֳ)�v��[6o %@ڿ�|�ԩ�'O��xl0ñzL�X^�c���<�L��m�|D�,�р�pL��@}t:=� 2|�!�'��b�=����=��QW�����B,���۽�	P3��ID]S2���oݾ�X0d��@�h`�`{���S�c��-�ͅ��|�g�Zg����ƉI���i
�3T���_"T�r���O�ǯ^v����{)��}�%o2��a�b�AZ�c�����'�V'�mq,W��b6G;�l~��-K"�8wAS����/��U�K�QM�GFJ��kk���թ��q�!pc��z�0�|��9�*tҔ�����d;-��!��_��ڶd�Xx2�Uwl/�w5C�0J�����i�!�r�j��"��N���*Pu�g��<�f�����3��O�?vbn�B����Q׏���8�4RT��W�Q)��1>ìiL$%�i���!����]!��oZRJ�[� �������qז���ܹ�3�ƪ"�Qő��]w�+�����<��P�����y�~qdxx/����sǎ~�/��C㋧O�>7pG�B��$1a^R �*��f� p���.<Q�
������s?+q�������dp���7��8-%\q�#x#�ò+�ae�,IԐ���0���m7<�`]�(<����E2"u��8b؂1�$���@��t$X*���
�Ѝb�얘:�DX��y�$5!1�	8�c,���y�� ��%���R�R��7����#����[< �z�� ���+Y/��K�ՠ�æ���"Urmgey9�ˢӵ,�r�'g��!t��^�C'�/�/y����a@י��6�}�	��5�>�\��L� ��"�"�Dš/��C��(8����w�H\0�/�zH>"�.6��[1�*�9�QzG��/����@C8��q��g+K��2���6���"o��F���g �����K��
�T�K�S�\���b�oKA���Ό= �`�P1��O�"�:���	FLl{�y/rn�f��X���P�u��$RJ�mG��`���Q%qr����Zd�6R8:�@��(.諸�{��1}��G��#ˈH@|��·=��i������Z*��a7T�fi"��Z�� �X�_ٗB{�)L$�(�$�Sr��h�����MEQ�їa�г"��#�"2~�[�=�le`PQtH��DA�t�B�C��W��z9tB�ci�T�P�J�.�Fd�$���Kn0�`k3l, A�xV"o��� 6��z�b	(�A���^�������tl:��,�EZ�F�Ju)��@w,�A�/�@k9:��Q��xU�4��s�t��H���5�h����[�NJ�2*�V�---�β%��T�b}>'MǭO*�/Sv����l6aS5��퇪�?<�¸땯ӄ	}�T/;�#�.�4�h�i�`�Aj��d��1��>�9==}�M7ѺA*�2:����P��!�[ �T�VJ�0��V��ٽ�7ްaUx�g3�DA�dPr�w9:��.8M�9r�k_��p�jL�Π��$$�	������[���թ���7��d��|���ؑ`�4�`=\��f�o��oo�������mw��/)q԰�=�o�F�|�����Çs��f�q��tQ���S�Z,�oߞ�gϜ9u��x�ȃ�i���.gux"�H�z�tX�3�B�WD!!�5'v�=ز�r�_���n��>�u�ʊX�����"�48�aM�Nc�&t� "��=�兑J�=���������������?}���{�O��*�빑�+�	$�F�X��22�H ���"1I�;�J�Ŀ/���J��1^�����MAH^�we]�5�./����8�̓ǎ�z�.)@m?�5��+OY�.l�^���t`�S��f��9v ;�A?Ӵp�0��f3!ƃ0XY(��V4l���ϙ����(<� �\:�χMR�eaKcLA$�-r�<R`*�����Im)+M��"��|1��	�U�:]�g� ú�O�m ��F�H�H�1L�!�(�����	�y�d�V�}	�#��oJ��=���l��͜<��Y�yVj��-v�l*�y�������fx]�&M�9D�Z��H�c��<���:����%}��9C��H`E�y�M�H�s'� ��Y��s!g5���X@�j���^&8�](�F%��t�������1�3J���tu����Rz���
=-���d��d�7  Gh@
(
6����N�ݬ� RY��(�I�2�{�=J+wp���aXR��&�G�>���+��#�Ȁ�=�n��:�r�����/.��ðbЏ�I�ٱb�,�����P����X�>i�FD�FК����'�k��xQ�dpu�o�G����jmqa��h"8��v3Y]V����rwc�,�FFF�?�8R�����h��.�h�C�M�`�
��ڴi�޽{�`�EpKK^�KDt��6���$T��b�`���B��:.;��V9D�$ȸ Z��	ʮ]�����_��a���>`��ٓ�D���.p
P ��a���gxԆ�g:p�gȪ�&c�\C����{��;����SSS�|�|�����ӧ�F)
8?NY."�3!%m���0�qN2��31Gt����u^�$�]��?96�cǮ|6F`MCڼA���kq���J��݃I�\�-,T�q��'Ϝi�۪"�8�	g²�ڷ�2�|��$9��^2���>8��0U��Bi�����}8�	{ю�E���{�����>x�ˬ�.KS14�O���D�t<���2��f\'\Y�.�/����C�	�&���X�8�( .��N��<|� �GӠ���o��e8#�{����+�*�**y�.�y�K8��Fw��U�ڀ����[!I����g;��ˀF��Z�����k�� t�֤�,2�o���6`�p��fa�UMI��"�B<�r����P5���*�K#ٲ�Q�������XI�JQ�`ڞ91V�7���i�az����<i΄�ξd閠sx�Zb�(8�w�Dw}sN*ξ�7Q\�K�o�~�!���d��B	��s�����~;�y�0�������_�cǎ.,,,�QEi�.�/��Js�pX�E �sؔa6�$\�d+�%�e��4���y���c�R�妢�I�|����曯;t���>k:^��S!W�I*Cչs_��$pQF D�#O�~�����g7v�����w�}��={6N��n�чRX��[Ė�Ȋ�d�3�n�s���h��0=U�{��&�RaϞ}����zt�R�4���A�C�1-Ca�������^PE1+��$�nD���lԚ�q���z�J6R�3;f�O�7�sn�s��A��J��c�W������Z�e�CHdIǎċ��u0�JF�#���8�gu�G{���ɑQ88p  `�|��ko:,fd�7y>vnv�Z[�d�l./U;����,Iks�oq�s/7M�R:W
Z2�ԁ���,%W&|�e�I��e1�R�Ov�|g(k�eᤎ���	N��R*��Ǥg։]L�'rl'�V�%�l>*�V�0F�Y�:6 �ss<@^��
�D�D
�]�ŧ��p����>U���w�N*v���2-��c����C	�2V�*	��@P,%��P6����x���N"�E<I��(� =& ݳ��/b"�m�!��s�(u�\)�jdi~y=B3��C���!���۵=+3�ٳ�k�%ǎI�1P9��F��J9��kp6!D�Qe��č-@.�Z�pS�=��pA��H����E�lИ�A�5�tb� 2`������w<�K���;�}�=�7mLYm���V�ה<�^�zm�2{xhI�BK��7:���O�� P6(��L.�/�P�Qђ�F%:�l\YR���fuy��[���Lx��%��F��1��q ���B(������؎�N����#g�0�˜�����Lcd��{vNMV���e�%K�'��lh�9����y�$*q�6�t34�NOi�lcM��i�a"J������6L����t���p��m�K".�J�z.�-�j���z��;��muZ���G�鄭�K��;۷or�C�t�� K�;؄��d`�bڤ��qH�~��$�#��H����K�=O�����z��Q��j��Jg�N��E%�׀�υ��N8A��(����w��Ȕ*$l�I� �X�����OD�s�v��hrrrt|��ނ�<u��s�6�x�	��� ��e�����q��a?4��1D.)�)ˈ+ᅖ�>�+и/��յ��ZM52��ܽk��k /&6l�vv}�:�a�A'7VE��z�n u���<�42�r⣏=��o�����{��d	m���?h�/��	�����t42����
>�R��W����pD0C�#�pu ��x� c�\����i�%�˙b�9�����b��� �499�Dn���tz%q���G��a�p";#�b� BwE	�I;��犕Je(� S�J�_9&��q�%g���R����0��2�IpU�~ǰ��}��_υ�uQSX���z�l���X�z�i���j�����{ [z�g�N'����Y�$u+G$%0L�����`lW��kזכ���)Wyf<f��1��;`��@	$��V+v�}����y����O�vٻԔ.���s�������>oz�W_�w�Վ��� Ӛ1 ~���f`�2���d 7�+�WA�k��&�j9sFw&=��a┉�0rnW�i* �AH�����-z���Z�5�ޜ>}GS�+�Fh0u2��>�^����� �BtH6?b�QX#̡C��p��0rG��� U���z��V��p��߳�Q�H�җ����~G4��-�%R v��੧��d�����#H�)4���>��sW^y%��$w����0C�V�Y�I��f�R���qLm��S�N` X�z�*�X�a���EP�	J��eQ2��1�cu<4,� W�V1f�u��ѣ��u4�T͓�X/�Z��o��R+���=|�o��7�vp�������g�K�V�����_������]�Z���й=�ۡ�Ov�Jq�^/��211	�4���	�Ϋ��
�ɑI��!$(0
K��M=���f�Mo}�S3�
�X�}	���TU��<� v��W�Ã=z��i��r~��=:m*T�֧c��j:`_�]�V�{=��I�^��^��?aw�<u�>�^��q���:����˫VJ~{����;���;1��{����~�~��ð����N�n�*t�M�bJ�pJ�܅�5~~�9$�el}�Q��������V_�}
?G��bQ�hA�I��FR�.:�B^�j��3W^~E�\�2�Y���
�+$	�s�t~em��Y:u�fZ�RJxgueݏ{��cA��ƌ�V/j�S������2ס~��U^]]��)=5=:@�N�f8�c;v�(�*qH$F��|���z�̹���Ϋ9Q�A���8��:� 0j�qK|���T�����u��9_ �w��I+��6�.�^���7��r���jh���H=�쥕%ݵUۜ�7z����m���.����a�����z���J�����qP�2�bxE��m��m��b�_9�T$T�K?�c�����"�Hl���=;���_����u��z�Npne���pԜ ���\Y=r���s˩n )6 ���݇�A�)��?y�T#����##������"C�r���o�dQL�%P�"� �-l-�؋�< Y���>]#;o�_�b�֏y��=p��q�0+�*+H@�G�Q?GT��K�"���c*o�jmlj�T���6>�y���m;�O�Lښ9�C$ ^��8�(�+�A�%�������OLn޲���)i�LJ*� �K�"�_�����g�~�qN.wq� (3,Sp����v�o���@� � �y���I�jh�K��f�Y�����ZA~���G5�s��A� %q������#��<y�% �
3�NL�>k��Z�e�yE�����W+Չ��ɩ���Y���m�ʨ�ĨB�|@OM�	��U�,%�%r�Ώ�H}��;{�����y�����Q�Rs�F��q�˕��e�>�>� ����.Q�V7��\�5v�qǟ������M3�4: ���cN)���D�H�ĉ ��RA�GA��R���)[�7���0M>��+U�����~!��N�_<��~�l، ���?�-�|�
>��R��2
jd��i�����.�7vQ�B\�4�eW��^�Z���qyF<
����%�p�G�k�����3�04`�Ro��w�L�5�@������l֣�B�.A�t$qI�Q(����q9�]�6��q�;�3��y�u�J�~�w
�����} �cǎ���؅���.4��G�%����GT`z�_QA%=��93����űDF�l� m6�p�p���u��R��Q� ����tj�wlҪ�=@��s�ioڴiy�����e׮]I�1S�ۄ\8aR�.��rB�F�����`6���4��-4��L�X,� �
�6��2e�Ά7����~��Ga�)�G�}��i��$XYY�����/>�����}���=��prr��5<X\���_y�d��)x�s��u6P���eXQ�ݻ������Ɓi�\[��-�3�2�K�lf�(��5�1��c�8q���ظq�{��ٽ7=������ѓ��N�6b�DY��9}R4x�1?����g�=y����lbygO1����v�a���c��Ϝ\Ym&�h��\�����?}�x�Q��Ot���3�&������\�-:�����q�Â�=�VR�l�ݶeC�QbJ�WT�H��0�ٺD�9��k++�0S_x�J��Y����R�u��+1�Z؊���8�5lr���gԲ�j����ҹ8��n���j��c'O����{]%ÄW�j'Js�i�v��������e+u�[�<x���/-�,a��P�G97�4h��B��?Nvr������S�B�1���{MN_����i��ǲKi�s5U�.�q�N����Ƀ'����?��>t��7�M� �AT�7WE�F�"�2ϵhm�#�ȑ#��������?��T����'��z0ʂ�9�+�e*��g������t���{��ͪ�����o��?���#%b�� �!��}����'>q�wRmK�gz�{~���������}��f�Yw������o�Q�� N�᏾�ohJޥ��O-n����CТ��>���=�Љ��8[u(�'-�O�2�P.��-�dS75��¤���5�{^��]'V��V�QӞ�����F5�䎒���?;�P�����
9/�^��1,�OE��'8̈́�}�u�ϕ��&�T�o�T�Be8�bź�`��M���Sōp�J�����C���6(�_~�����驑ƨh��Z�k�jcz��sX�U!l&G�2)����[$N�|�J�*�݉�<�U��g����BU�#C���T�O7�����U �US�r�
�F��(�vK��V��u7�깵#-/.=�P)�bV�[6��3�r�-�fy��8V�v��4}K7g6��l�5m:�^u�1J�JX�
��%\Y�p��}��׉�.����v�� +����|+V���!������;%�ڠ�*u�t9��n�Хr��2S��LNn��#���]vYmd�k}R �иPpjK�8�-,LfjH��P�9�	u�ǯ����9���������[u˥=�Z�kMc}b���)�x�
��L�|�h"4�P�rmrvn˖m�3�F��
�����9D��N�P:&#!���d�;Gv��m޴uvf�^�A�Pȫ�-�ԍ�R�,b�\��4Ŏ�C?��96L�N��ݡ��,j4Fv��}��7m���5#&g����&
�����Õ��}��7��<R��/&cX#����~�UW\������o��:������s	�j;7�h蒌�O�T���D�16�ږ���N�\	3(%W��Y���ݴTn����i��pS�ajf��,�z�^����\:��������u��5� 0c�&�]�������PtNu0��W�������k�yW��a��l|����Ï#�a*30����6���8#��Y��?�e�T�k��c�
��",�@b%�T*�h4j�,�<91}������"�K��d<��v�D�x�����9+s����̟�]�t7�	QغB�El�娗ns�>_g.����h1m����)<���H�G��HsJ�*b�O�*K�T�-'��.���utt��
8S@��/I	��l�IC����X��0�ĺ��H�v�s�$+�H���5���|�qb���P�(+�O��i��I�o�}���{x�� �Z��g�X<w������H�~��i�8H�V�`)�R���.�4�D'�od�Y�K��+5|��ɳ���7�p��?zt�������G����v�ܹszzr���+K˔iX
��C�Lk�ֹŕ���K�����Ť����p]7�>l�9��s�9v��^i5�۷n�ᆛ��8w��	ؐ"割ɥ�Բ�Ն"���ӓR�5,���ɉ�ɩ�Y剢�љ7*em*LN�QD;����4�]�911FnJ���)^x�
��{�گ�['̎������N�A@}d�+�g��R��\ĝ�ߡ�n�Y�YidX�����������b[^�ֈb�eQ&��2�u�A	�b]a��x�KR�d���.��ܥO�6��t �?� �l`](��/?� �r���.v]��Q��̱�V�xݕ�y��Ni2M��q�F�D�9���7�u�=����y�2�y��>��?�ɋ/�t���>�Xԣ�_j�A��x�Ǌ�w?2M��o����o��n����=WlZ�822��o~{u}�4��"f�����O}�C����=�v�2��Ywサu�N|�V)��o��~����_��\\������ﮯ� [�A�X���7^��_�x����A�^9v���Ԕ�w���Ƒ�D��>ی��a�;���J�𔨡xu�<�i�$�kv�FJ��m#$���8#6e굣9e�֩�V�Q܋�zs�
f޷�
�N�Wo��9�1t�EED>h�*�v�UGF�eΪ�'�$z�Ʀ�6,̻�2 �W��ϖK�ͥ#��<��c;�f6F\�hS�xS�,s,�$��ҵ�U��n�ͮSшТ�h��2%�'��ļ����`;�r�J���Hz=ᬜ�|3'[�nl�� �Uw���k���ؑ��O��ᅰ6,st���H�	H�o���kk���U@��[�LOO��):�;Iv��4'ӎ蛅R$����9��!T�iG5)[o61���q��#k5����}ө�u�l�l�C�+,��9���ۡ�[�E�\���."��hq&
����@^7WWY+si�-~0C�2�>�S�N�[�i��&�Ѡ�NJ��"�D)�D�F�NĶ�J�M�5�r���]��ڽZ}�?R���n$!Z���6mh@��)1��l&(oꞬU��>�5�\yY.{Է��$@qWma�P�%�92:9%��� ��2�1R���k�I!�B5�o�,��b�$�D��Q��sff��m����`W�&�B��v����o
���UBZ����OcK��m�7F��s����z���>���ns5:4�D?g�AF���Q09�6j=`�"�F��q�5O�)��kl��	�ES��4�ņ��!H1sԐ�����tI��sOpm	Vp$bªY����R\$Qg����_^Q��;��'b?A7c�98�x:])���[Q�=��4��ᏽ��bj㌙ͱ�+�g8tPdJW�HD�2gsq���V)s2�;�T�OS�5����t��P��Q�|�-m���R����`\q��S�p���E�s��0p`>n��"S�x��Z�v{"�D��0� �lj}��#:�������膫e�CF�Jy��m�!05�� �G!�Da<��.0C�|\	�`��#C���[%A�F��)���I�y��^�p���-�!���*ƒ!2��Ab�O頇R��NdP���ɡ�51&���9s��ò�)[S\P�S'{s�"�5����W�V[Y�ٳ�g��^a�Q����k�:U7��n��?YN���/�+C\�3�l�(�!�p\#+ҧ�~���_]��􉧞>�ꡍ���������!�G�ƝS�]�8s��up� 
k^�\pj�(�\�:Z�=��������?�i����?K�W�&���$�6�O����4 cӰ�4����q��u�M��®%�!�2	#`�N>HM�lA��k\{��ڽ������˔"(�B��PG�F9��II��sDW����k'���[h& @�Az��{A�	��!�(�$�@�Q�fs-摈^��CJ�
� ���A����+W�~Bc�A(b���ݕ�ϰ!4!�XШ�	D�����QٟGz���"���IU�&�,~󘻃���NU$s_�̥�J���D>�S���B�Ff(G+�%������R��M�kC��F��g������_x�K_��/<���]۷*DeUP <���g(��5e6}�GU�x�;�����S7�r�둺��V.�t�͊�tb����u�3��]{~�c?�=�a�&��c���c������c��g��.y�чl���V�ŖaO����G�k+Y�b����7��GM��6l� *Ă�,&B�?9��Sm���$��k���
K�{E�C���Q�~��tt�j�ˮ�Gz�GA�CC��)>�Doм8U�"��e�����u7߰eF����=��݌hF�4�1�����N
�%�K�A��n�t���٦��Ǿ�����pU�-t���U�Q���T���O?���|뻎7때˶m��8F���*̅2��Cݸ��&��⇩`QF��Q�ݐ��,� ��PoP:?�Y��^~ͳ�"�S�bGlݼ!-��T�w*�T�Ӏ�bQ����p�$�V�D:\�Me8@6�cny�لu\w|j:Cc�"ꭵ��k�B릚��j6[�lP�1n*������r�: 4kk�l�u}9�u�1�v�	S���)ԥ+��ԊA�i�m�t����#R32cJ�S�-*���Ȩ��N�G>)<���������;$�jA��D��8띪��uDRJ?e�m�Z����u�ݜ��n��NM_l."'6�Wk)Ь�X�^�y���Τ���u��q�*ǂ*�K��pچ>eu{2��T�0?��*Z]��ف
l��p��>1^Q~��MK�T�j�(��
;�F2Mv�(������nou�]�Q��~.���������ԅIe�4v5�{�*����^�;���$X����zٙD�h�"������ c�W�6T��iu���̙s�w��]���ھ}��=��G�豓g��C�����i�%J㈊Q Bl�4�&�r��C�uaN��7n$l�X����
V�#D^H=>
U�w���Aq	
!|xuyx����4��L0�{�"w���(W�z)��a�Q��m�4WȤ��$�.�'��"�`��a(� ��׫�~��^Ǟ���2���H��%�"F�Dg2@0x�ӧO{��=Q�UY���^T�eY���W
��Uq=��Zqg�6� d�89{�d@��L�����_�L<�����F�0��E�_A/c�b-_[_D��rm��<����>�)�;���EgYy�@s��踅����BƙOZ�ُ�X+TӶ\�N��"��W6ء�M�
ȷ`f�z���S�N�bc��x&e���΋,y���Ѽȼb�
�`"J~e����I%� ɨ�YnpD�q��������%m����aa��o�-|�@��JU5T����s�=s:��}�u���.�&��8�-A�p"O
�
�r4L�jioP7H}#
�R�]ZZ������\�7F��C����cGmߺirnַ�c��:T�a���06���:$A��Xݡ���N���:v���U��#ľp���g�~��k�-U��g"��tڞ�%�J�4�g�9)gަ�C,�̓6l�z_�22(rJLQ�� �nT��J�r+����O��ȋ�vtj���VS�zxt?Ot���,��iy~��a�JT=NٴJ�4����Y��Z��nZ(�s�E�(*勳��-"�(̡��vU)7O9:V� Hz�T�	5>��ኤ���Q�<� �R�q1́���Ey�C�R��А'���j�Ի~,H��x�3�*�^�� �p�Rb⤍�f�Z�ش>dy:����/����O-�=	C�J��E��=|���WS���*���0l�B�%׍H(E����}q�'5�A A��������-�ޞ��M2�4<���|�Ý����/�k�R���9�m^���'��w�]��+���//���w��ΡïnlL�j�[�z˶=���W.ծ���[o����V��@�S�l��>���폺k��;�+ui�V�*칐�q������gA)ۦ����F�Bp8��B�;���'�(!{��0� O�j�;�`&�t��*;2�"2�f��3Y���-��o~���~�3����-��S�r���rK1���I������n�8:�3�4&&�ƭ��Ž��;~�>��K��2���/L�E��Qb�R��51���ijo޴kfv��])ʅ�R�^�^2t��mP �©�[h�HhJ��`��&�^����B��9��U�I@���g$���׽�ǝ�X�r	�H�r:����P�����L$�ψ� ��peۘ�L�;�nl��[e�˓���ky��F�]T��^�0pao+�P3��|�C$;*�["��JT���@�y�"y~GFF����(V�Z�sc�R���`D�6�z
�Ȯ,�W���Ř �-���B$�L2K�>�b���`Wt��S�^pV
KFMu�>1�)�!�QSɳX��Q�C���Bbb��\���CO�i1r�j�h��c_�P#�b.o�i�r���Z���V1ґ��}����L6&rN\��i*8����s\�_�U�!%�����*�P���^������?�4��o��i��*�W��4���̪�}���"`G�HaS4�6�N�!QS����c�e����_<{��~[��G���AųK��B�va/�%���@89�n��� P�ٵ�����q������|n�t������E�kktZU�P��𞉉�'��"�\E�p����TC3��WJH��\"��<�������w�'�<�xF8U3˦N�"F�����o�����[vP�e�i,7�A����HO����@(��̰���Gl'�	��o��^1l�H��K��c��_b�a\r8?D,)�K,���2� ������mw;�t��'K/pCgY D���&�ӄ8 ��
>�<��2�d)˺�5H@�b�͛jͨ�+"lb^2�}�ۡr2�2hbbF #�6�X������+�,%�ŷ��J[��c8���|ʆ!���eV�)���\8��p�!�C��<c�Da�vyS��;ur�Z��N��)5mllbTUl����<w�j�	�D\E��8�;�j�}7@���
�Ԅ�/D(����s�[)׏;���)q��j�Z�u��g.-�[[Yްy��ie�
���ۀlI��(�}Hu#��^�F9�U+U{D�s>��<�L�j��S�oU����V�4D�r�<�����"_�/乩�㖢�c*b�Vr'הH�=�{�Qs�����قM�׻'O�ܶ}���{��Ɂ�;~�H�l�٫6��a��ݾP3&8l�(�� �=����(X%� ��u�J^�g�����Y"�@�@���V�"ڍ+B	�f��t��:a9v��������-|Ų���96��3]��%sph��r Q�t���P�MGU����<�n�K��z���
 r��e�hrʻ��kv��r�~�]q�c#㰡�w��@���WK�5>��fl�v|?4tj�1)r�ω�T7���Zs�'E��I�gL��ᥜ8{����לV��{�$��~��_~�OVVW\ۢ><�YsR���tT!��Uq�°��O�"%j+bZ�Tv9�W�VJ�"K�0p�[�������o�=Sl�@P��]ز�՜)�r��m7W���_���o�����$�o�������t�ȋ�5P
�K��}����;����=8��S˫�Uk��9%�q.ku*b��K���-�`J�)�j��M�n�<����<%��Z�a��Җd	�$S��,��h�5��Pp�?Ir��[�	�=���%_V��]�J� �5R�k�3�3a��|��˶)I�	U�k	��$�rYeD�2�uh@"�Q��w�o����u�C_�	��F�Q���ff'ף����m�v�W�� ��P���}�7W��!"�K�ΦM�(=�P�0߼eK&��@���2�� a�î���&�c`7���ժ#��� 2�{w��&��V�S��j��9�'���&)�5��.�"5���Ms��5̳�2�����|�D{��5���a�$��j\��D_?f��6UŋDd��0�\�f�ԣ2$YL�P��`��ס�ų�W&�g+�<��;99	X4�f�I�����eU�u�)Ĩ�cIT]�}���L���,�aSXM|k��m��T�taSI�F��e|�'���)��?�� ���b~F���[w1�jfF�Đ�7l��˸�3��\���Ȭ(I*�K>��ukTH5�.�XT 	�~Fx^$�4;������8�,#�zN�4�ANk�
���ꗅ���<�I�k�.��M|KG����kKd ;��Y������,-uu��(�3��{�������bKXz����.�o�=?ڼi˻�~/��~ojf���\=L�lY���JJ��*tS
84L��z�.l���<1�i�r~�(m6WWW������%�U/WA:&(���=�KD�w��pPx�Iҿ~�f8�MYs�@��C����B
� �p�?�)i*�t�D���"�$�~D"f�FC��(�VI2n��d$MNŰ���4�$0��W.]V��t
���J?[�M�z$�W���v��nO�a��̾�V�,�	� ��6�lS��_^JY�q	�����EV�\��^��Z&��[��v_@���h:r���}J�BpsuJJmy��;�6Q�0 {FG��8苫q�Jӕ��s�@zg*ע�c������s(C�*H�$U2#��a�I1N�9�2��J��
3'��zM�u�%B�q��µm0ܒ0V��G���2xK�$�����ڼy�R��������AI���1Q�������*��=e�]9����}p�����1w�ބ~�� R2(�)�d%�"�j�T�v��@���X&&��˶�r�-��(F���Y���0C�3s��l�YLS+���´���1<T���_`��?I��'������Z@�A&I�j��qfr�����x���9�aK�;E���+o�&�+���ƌ)Պ'܂@�@}��@~C/�sSx�s�r�R���ۥH|EеQK.��l���+�_��C�8�kK����A�<�Ƙ��1�h­ȺA�e���	��("tἋ�4mT���#�^{�e�|?^<����~��_�����o�Χn��v�Ѓ$ܵ{�����Ԥ Z"�D
���`ee����a;��"���v��{��.���;����߱0��F~~A�N�^��ҝ0�˥�^����ؾ犩��N*r�7�!�BSN��(���A4�Rf@IC��Bf!�J_�IO��W�Z(o�2!�M&&��}h���,	 $�V/�F�Z)4%�z��C���d@8$����ru���Ĩ�\���z~�܉�{�i�, \=�י�^���kgf���r�jl�z�BaRK��x�)����k���X��ǌN[�AX}��2�=8ï��%��y�>C����NC�Q�2�i[&�7�h�+W��H������=�M����u��7} ��p��̃b(l�ߴ��k"l\�6:�\�~*� �� ��9|e{�&���F��������Oܨ� @迟Z3�q�B�����6>F����c�6ur�a�[��_�?�4b���ПظR�_���`FM��3�Ҩݎ07-�J�?6���U��x�_ɬPrB^��y�s�M��.���E�H��� H��]�(W�bl�$@6��M�R������h��h�Z��
��$MZ�M�l���[���_�4;�������E[�hxezrbm����x�퇉�8�u�4Y?��Z�w�����j��ˢ,G�&��U��	�ZW3:y�%ױ�`nb�0�Їa#H[c8�bCV+PW�=��Ï?���;c���������jU��2�(B�*Q�F�e�J�/�?��˯,.��Q��!�"JYOS_��d�d8C�����H�Cv"�HƓ��m\�QDh-i��ӁT+�?�5Ќ�˖�3�vF�p���D��Ydl���8d�E}Bަ�)d<�y6R�֓�.|"ب��UL�d��	��<%�駘Ƒ�j2琚Q���u�d�@�%���Xcg>	�H!}Ѷ�_/aJ��S�)��~��?Q��i��y�V:���r�e�X��x�z���!�,��V��Q�j��P�
6'�Z-���;EQ�gL&�o�>X)|$A�Ǩ�����+��˫���ַ�{�9`�Z�z��׿��;���>��!�(9i�fPJ�0�u�j� Px��'G'o}�VV���*�y�u��p�M�6�᮵;_��WN�9��Pa	[ҡ��I�re����A�����0M+n)��a"~�[�B����]��J�g��m������{m<~W��� ��,w\�Lt��8-������!35�	/v���q�KB�C$k�!sBt�!*�Q���w��}�_�������d��Y��@���.J�c�TGA�9��%�z^P�C�R��kIR���hI���k�6����y|�u+�W��VW�?�ן�{�{�}���,D�m�(]���䆢���jUO2����ĹX	��\��*J��A�J� ���y���R�*����ݴi��~��ٳJ�J�DrH�Q%~�Z�2������
��Ձ�m��R\8�z"��7o��|�����d���������Ϟ:u���j������ozӛM������;�Ϟ�}G�CP5�^i�Msf����Fi �wvq�o�������Cv
C:�n�Q*Ta��R�ᴾފ�D�)�}���s/=��3��]^�>/~ �)2� ����.�r���!���7�E'&���G�8�`+X�"��"��\ޖ�d�4"�g|��Ĩ�i�+������E}�Qmj�Cnȥ�
���^��;�X� |T@��qW�ג��$A��ǈ=թ,�$�ƍ��p���G�\�ku�ؕ�g���aS�^S溩���Z82��S86�W�^.sC	v��K��Ty)�w�څ��e�˄���ŉa�$�;���r�~ƚh.�ͯ�Lyr���v� ���u���C&�ev�B�s?'�s�X����b��k}e��W6S9�H^�^%�τ��s�;�!��'9�O>)��
nB<�HR��1|�u>y��!hL#���Ѭ��c��
�����]�!
���[̩���h���O2�"��0��B\rc||�jz=N�ǟΝ;W�Vh#`�]��c�Xk&��E� ��|3��a��YDď��k�(���2��0��oqދ��aZ�-|��<N����W�Ç��$~����3b����4?#��wfgg�p�]){n�[<�cӻx���W_}Ӎ�S�LH�x��鑱'�����ѣG1��Q4�ꋧ�R:���3�Ɓ��b&�����a��A���v:T���b����6����߂V�$U��#ēb6V����KQ��d�k����q�Ibb�����0	��������/|�r����vWĶ�d�8�)jb��m��:~'KG&��4�����?��A��?#�[6\�R�8wݰ[j/�7�C�y�!u�R9��E���3�Ý�u)���K9��,s��G��b�+Ud
(M�~���
W�0�{��u��D�kM��e�G�l��|{a��`|e�I(Y��:�˶�#��'���8�r2>6�\�pY��`��k�
�����h��Q�,�v��'\���Sǒ��K���� "�v�ZZg,�l���y��^owt����\�Ps���P-�lj�f��b>�Lp����v�p�@�ܹ��~���~���S�N��RI7�zۭ��ٳǫ֖��VWW{��I�-�<KD(��%|"��lh�];7��-w �?��C�Ν����[o��f�0p�����%qZ���f�Rm�["�BHЦvm=�2�"�scN�,<�&ڏr	��s�?u�!�W�S�HY-�3�@��9���Cb��lo�0�Flve�\�t�2�Lz@�#�wI�!#BC��Bt��.u %L�%��Ԩ�n��_��z]�v(ڦ䪮�n�-���z��jՊv���� [�4�z�<h0Z��^I)1íFlO4��ȸ7��	��3��O�<�=��t���3��l���T�DU�U�FP����x�M���=���GFk�f�Q���q۱���ǳ#Ƚ���t�Gj�0�Ο[�;�x�0335??o�N�\o��Lƅ��]Ai+�����E�t�Cf�1��c?Rt�ȁ���
('��qp��}�Q�];w��&���ӰUՂ��y��o��'��o���Y�q�ͮ�?~����/�������K���z�[�c��t�[�U%���v6*4��g��J���>T.�x:F�|���	�v��:󹄘G:�~J���fW8ӰH��K���g�FCU���������?���R0I�х߽�Y�AL�bOA�}������Z�4��e�J ���Z����pj�.�e�ZwM����J��A��Ć��i�bt����ַ��~'��̙3�������/>���ȼW���]�E�%�60��Çq���۷cǎW:y�$̌��a�MD7�������!�aG�Qi���B�`3;v�_ܠC��.N�:���Ô� ~N�8�!�!$��r�e�AO`��}|�b�� g�D=C�m(B��h4�>;VP��XVz��l�a����&fC��`/���<r���-�^|eӦM��0'��#��^�=<,f ���$����f���cT�J���/j��q;p0w�'1��cAfyb��[`-`���8��(�n�[�l��0'�4\�R���Qḩ ]�!Qs�o�Q%����oJ^S�?/�Bf�9'D%�g���w��1��]ۉe��h�܌t����?�)&C1Y�Ͷ�,����V�"�D�y���eŝ7�:��K/���^s�5XA�<*�V��Ҽ��p,��~�����*]1�u�����+�xN㔚/��J��U)�%չ��E9Ry>:RoԪ��i{N�u*iF&w����o�8>V�u�gN������N�Yt�҆�9V�6�S�8�˭�:-D�Z��`_aM����v��β���
Meʂ+�>Y�����Z�8�U8��<ܦ���Mmt|�TN�@7�E��Töt�hv�� ߢ\��1�F2n�c��N��	��!�n�&��,�z��Q��8�pC��N��;�v��d�\?����
u��� �(D�_���*�T�E˹XJp�0�/�cY�n�B���d̔����Ik��x���d���$(TM��0�o\ɂF��տ�')ߨ�$3pq����Z�����I�u ^77U���t.�ȕ~��~���&���V�EU8���޲y���JѶj������.b�3��u�H�~!&��Æj�#Ȏ5��_��?�S�瓧OMON�ʯ||fff����f���u�C ���E���\$��+��tRz��#������
�u����o�k�^=(ڎ'g�V�\vﾢ�my�Ur]J��{��ZԤ��R-y��㛶N}��5f�1N]�9�t��zE������(\�P��.ɟ�i�8@�����
�_f��52�ɵH��x�8/��'i�P��^�c�A�Q����"�Tf&����Z��iN�^n��ь�r�Jc����{�f�j||�*T�x}�4>S&B-�~���څ-%Q���cB�a�t����	��w��N`{��Ԟ}��>�׏=�P���VV���jV�7)M�7�Ԕ}dl��N�7�ۅT#Cht�V$V���j�a{vn��G>|�u7�"ԝ,�s�r�rQ/�y�5czf�=�y�5W\D���Ϝ��w����~#�z�� ��>�
�`Q�4R��
��b�/.Ԓ����]��m������9(�'����a��*�^��=�r���W|Ϋ����w��6���?�3����cGO,5װ. ��_}���{�ȑC	g�t�-eX�g�~����]]\2Jf�ܩ�0�n���Z�j³p�n�H���Js���O� fe�Gy���JS��ۖ�
�a#EB�	!nhI����7���'�N�a���U/���Ѻ��G�]]ZU����i�[\q�Z�آ*1ʫ�~bYP)%���`�$8]������E����n�Sr�X�-�.�T��N��ڽ���w�s"����1@��G�3�ğ�����\��+G�R.�x~I���9��~��g�ڮK�p����%�f��>Z��V�759�w�@�;�O���1(x߽{7����W��''����͛�6�j�-6[�1
%���0
l���qA�
�����O_� �`�[ŗp_n$�K�WذL����e<�������<��n��Aq��m�6L��#G�{��xf� pz�� �ω:��I`Y�a�T��*7n\���y�$f����4[m,0=�E�
���z
OA�Z���r����ټ6���f9���}�0^~�e�W��}啃�T�òb���Z-�ű�r�"�S�<oVW�a����Zƃa��d3H�kHd��
&W\c#Rq��A$'��f���"&��� �-T-3���,/�&��fY���,�={���0��ZY^����@��v���z��+��׏:r�8٢��%9�Ѹ�T{Ќb`����M�g�At����������U=�i��b�T��/~�=������c���e ![؍3SS������n�l]8���܁���?����<�)����uJ9VI�g�B��`Y�,K�g5]ٴq��j�NM�qhz���Wr؉� �4"�2Ѷ��^�aJٔ�[�,�~�U������p˿��qT(C^����x�3GG9�Ħ��ùʦJy�����p����C-U�z=Q�F�h����x�(�^-���qS��&Z���?��-ti��Q�~^���+�6�v2��R�Iz��ky!�l( /� k-�j,��(�h@��d:�Q�޽�BIF�.i@)��5B2g~�FHڄL�"��r+�֘�����"�T����e��?����'��ٵo�US���j���g
��C��O�hzzz�޽O<�S��X�q�i�=���Vs|tl�ƍǏ�����R�2�0�?}T���Tt^���l�B��@C�wu�*v	�
U~4<l�qد��5���s��O~�:P��w���񉩯��W8� :�/=��N�ڴ���8�����~��>�Q�rQ4�k)D�~s�]��,!���r�Nɔr�Á���܈�%��5��o��]�ǩtl��{bO̤*}��p
bQ�EE�
S��S6_�IۙH�/R|+皩�j �\<������/?��#�V��aZ��(�u������hlls+�Ŵ���������<;5R��2閍��z��}���Q�^��S�iw��8ѻ���~��'#�ZF��[ojxU���̙i���Й+�c]%���QR�5�z�<���mmݲ�6:g������9Y2���UJ�F��4;�fj�T�w�ܽ�
������=�PNWdȊ��(
���(��^X%'���w���5	�G^���DɈ=�Zv�P�V-U?�ȧ?�i��ko�{��i���FG���'>�����W�r��a�v9n�1pl�֘��&�ra��E	a|��J#��5�R�u�:]�Q���S��IsAJ
�X���ܤhR��LŶP�z���JK�<{�ZA}�R���>T���.��j�9��ѯ��U�օ������z{*��W6S�{A��8�E�d���j�kJ�-��6~��]G�<�tJ%7
�dBj��C�N��q�)�ڜ43&K��G�2F�\ ,�k��3�����=��裏��X\n���c�^�,x�	+��Z�i�ũbڥ��г�+�:35��2/�U��a7�m&��*c#�k+�YB�/�@�0G�Fegw��f�3��"��G��S����QK�B��7��Z�-�9l���b�Æ���\n� ㍕=fj �2!�R�r�����,f���x����i�e-�C��R���iѳ2#���;�.p{������#4]������q���w�9p� L۴�(����k\+���b����FB`�˾d��(Q�=��P�"��g<�Ar�d�E�@��R�}�#WƸ��tqvQf?2��^��V����Z�t##UNzd?f`#�{b��}�"s<�Vm�D�$��C�ݮ��\���	�	�~�ȱZ��{��Z�,�#�ѭ�ZH��*R�O�M�K.�Z��=�������Rubz�^o��晧O�8(�e�浵�n����`~a~��z��i�2�7��u��G!Ehr�fqRp���K�)-y@؞Ѽ�ҵnkuy��e�7�*upЈREz� ��S���$��>�ñ#GϞ>C8$�5%ު�ؐ�^��5�$�fF�E-�fL]~��XDCWMM����L9rq�-}��Y�c,2[�t���y8iF?PƆ�6�T�U�Ҁa+e8�L^J�e�O��u-O�	�eY?�M�A_23(�y,�\^�#BJ�_h�Î�)�䶖�k��o��l���!-%~:�θ�+/'d8�k���g'q�m9�h|$9�β�����}���;GL=�U;q��c�=�u��+��w�;��r�r�����2�'�"�dyl�g~�7����!�GF�r���D��
���������<����Z��B�k�[�*i.2�,\�8
��3B-�ن����R>����m�7�ϙDK�;�f@Y�K+k���o�U�� �R��Z1��K�S��-9@X��Ҿݛo��f�Z�=˭��݅J!.%�'�@�;JJg�e[�{ ׎9|���0�-���#�LU�bDVq{�#eg�L�d�~Lv��]l�6��9����[�2-�=�;���,��������g^|����'�~��)���R�U@�Bpf�Q,��u���c�|�E�f��)�z�������>tχ�V�J�P!(Yd��Uk�bDY�xU���\�в8�)�i	rB�]���B67��ͷ\�T�Y�ۖl����;~������al���Z��G���������� ��5�-�q�����^�s���'�|�W^���(�8N��}Ѿ�)Ϝ3~f�}7;�o,�q�=˺A�^�U��\�)ըb���)�̩E�f�7�1E8l��}�������U����J�eA�( P�0l,�ܽg�G>�a,��}�8ǚj��(yt0{]��ܐ��#��f"
�K�w���3\w��3���I�统&���@���������/�.$ĠD̰oP[(g�.����@7����O��?k����O~�ڽ��W�{�P�P�8��"%�\�c[�Tv�ں-((S���S2��5��*�6�[@�.?v����޽7��-�Uj����&�_�^��+E:�-��9=y�d�R��#̜Z�g�u�w��2�5[���\�a}����RNK��U�7�י���M !��I��<�=g4`��0������(-����*`�l�:3���PN��v�葅���s��i���
Eáܑ�:�]���± FN��Q����:\��a;v��8ې�s��|�+�9.��q��q�X������b=�Z�1(�	%�����Kw�O��K����O������K/��9x<�l�=��s�3S%�YI��$�5.��tLl��
X>��w�{���'/3)1��0���9��}8�����
Ot��Y�$a�����g��ѮKa@F�!O��T��Ξ=����4ɀ���ֈi;���zs���w��&;��Q�w�\@?�%˙�h�*���s{��w��B?H���A��u*�B�P�]4�k�Z��0u�&�C�4�{�W���o�~�[��N�Џl���l��r���������oz�	_Zm2
�TO�{6�%�l����|���=�)a)�(ZZ\���3f'q�j6M�U
5#lW����^���u�=���OfA�V����;r�N�'7���X~���tmR{��w�x�-��G� ��,y��G����D4V"��Ų"lԒ����5fD�("<���Q�0p̊�KT%T5�bcKSGf屃O��%w��$p(���*8�ӡ�_R�$�z��pn��Z�(�c�2�N\���R�����U!ZV��McAwɖ�Ħ|�٪����KE��.����� ��L��E���9�U^��X����n�Z�&{�\Ro���,ۂ��Ǯ���w���ڴݔ�}.]�9[ݢ(3��"ވ�k������>�S)���;B�a���\a�n����DΠp­�b`� .���|N��S!?� R(M̆x،6���(��ʵ$g��q���ko��ٳ�>M��6�`����kD��{�j;�Z���E�uG�8�F܉k�E�<6��/�Ls^$�f�:��䓏�>s��s"��Y��H���[�(�Ԣ�"�lͮ�u������
�5�k��R&���� �DcMXf	N�M�bGPʞ����4� o�����Xi�IshQ��U�����o{���4�X)׏9y�����3a��2$�C?�k���.��@�T+�8���^�-��|��()ZѭLWG�#�����R��t�㚍���?�}{�����T;��{��_���]q�G�js�2�_x6����2�v��E?@�� ~vy��R�ث/����[\�A��ɗ^>t��Y�W�iW�p^�r��@xO���P%�|�w�Ɉe������<��K�(�t/O�#G_��ګ����������G�f�<� �mo�m�e��Q\l�ڴqn~�慲�4�۷�R�u?h�+�����nw[������^P�+�w\�p��W��M�i�n����+.W�rA_k�\���B�C:�1j�)�hBVk��"�棣���0t�ێ�$�J9�-�6�$ڢ��<����7nPH�����3�������6���X�]3S��Tr#��0���D�"ji:�
��$5</섭�V��X���zXED�[$��A�^m�3uZ�4��Zk-_���qǅM���uaHj�1:52 W%���"�ә3瀺F��M����aW&��hǎ� ����Y+�g�y#.��F'��R!����� ��(��tYش��k��{5
'Bˈ�'���Ǐ�=53N��N�M]��0�\����c?99�4�|ʗ��W��͸�7Q�b���{hr�I�Ն��@Fޜ�ŅL�Dez���q�S�n�.R�5O�Y�Pk92y��C�Z��q�f���je���9�7�>�"f�����&�LG4�^/�T��C��[^^�6��@�ںj���՗e��_��F'�q٥Օ8�-�m�OPg'�ݏ�ī�L�4oV���c\��a��k⹘O�����1��8������)I��
�e�l�p1'�a��x���5�b�
k�c}���alHI,��jc�ةL#4�(L��:�%&3M�r�s\�Cp0x0��p"��-E�"#��b[����,�o2M�nbj�w"<��A��+�\u�n|,��$ ���I��e��-<ޭ�k붍�Μ>s�혮c\�g����+�W�x�T)?�]�|۶m_�F���3sLŜ��m�ˎ�����,�a���@ĶVWE;)cf���̙��nT���tU-%W���	H�j�� #�M5��j�Zo�����?|&l&۷oW-`n2��'q�,���x�)v���/�첵��/�t�C��q�Y�I?\�u	�)�q�rÆ�o��޽WF��֨�>�is���m\�u-��AҁڿR�\���p�)��,�OƋ�z�\�{�(�a�f���YEi�Fr���~����8W�$I$sHd{.���+�}:�1B��pGIh.�B6tMm�8����F�5MD�Lpd)�c�SF��n���T� ��%mr��@2u�YD�,bߍ,�b�|��;æ����+�Zt�.!{���E\��盉��4/�5�m̲����45�g�4Ujel���i��[�n}�{޽{�NײM�$h09ٷuU�፨-	�Dy�R�ۂ}GY>���;<���P�C���Ker8�{�k�񉩙�M/��r�w�o\�"_)Dʟ�..-�Q�c?�q"8i�#�&U�Qb�R�,0C�ul*�)2�Rlǫ׫�ϝ���e�@�$���h���^�xQ�AiT��S��(�Bp����dF*x�H���)g�<҂Y4��v�����3����������Zf���eb��I�)Ӆ����HB��"��س�q� U�W1���	f�bEUR�~��b����CZ���vר�HJl4�n��o�⪒U�IJW�l���L��;ݚ��N:�f躍�����	qw�Z865����;�0�����c����o��)�s�,m�]:�����v�͔Z��T��)Q���w�Z��J��חE�y次R��4��۵��w���ko1m���1a���e�N:G��ꕬ��_��ϙ�=n��^��Z����<4_�����D*mXIfc	��-h`1F��{������t�iQl��5�K���iu�3 ΫE.A����,���N����ڦ���!u?�_Z�>����/�>�D��J�}���7/�]=vK�U׫���6������_��3/���3���S�z����������j�[�O��_y�A]��Q�\������S����{��z��a��[����/�����\}G����H�ƃ��\�K����!Ĭ;24D9!�(ƣ�B��9��~'�VA!�"a1�V�C��o`���N�� MӴ����KͬP����w��օM�a���:�kg�ըT�Zv�Z��<�]�Y���׀�K�n'��"\*NG!�=_(�\P�xnI��N8T�j6�;v������f����|� ��ܽg�%gv&��f��Uu�Ww��ix`f0��Y��	�2Rh%m��� J�@��bH��rcE#���gH��@��h����]޴:�}�=�����@�P]uo�7�5�y�y-0�Et`�X��tC�?�!�T���O0��D���idb�:�K5g�TR�[��z��M���O��G�Y����W�⑄7�E��ܑ:4)FQ��P�Bפ�H�B�)Y}�O�!n�@�[���"���]@6���~�fd|A��>N�ʠw�?�A��S��Bv|T�VANMoܸA�幨T��4x��#�CD�j��4w\�r�a��'OҀ�g��P�h�Tf���r� �h��z���������T�i%�}�TuS�7r��_Q8���O��scSϓ~��TaG1 1�Ȫ�Z^F� ��GH_$�G)ױ@z�.���PQ�f�Tyq:���B��p��$~�z�驀̐n���#Fõ������������\M�ǨW��>({O� w|�X�\������{w���򫿶4������4_({E�ۘp۵?�O�����.1�cǏA��Ν;�/Z!�9Ys"�z}b�-l����YX.�Fv?��&�[��'#�*4��q,���3s���澩��n_m4���l��Q�a*���ں����?�������Ugg%�O��G���{4Q�jIa�Ѽ<��ë��yC��Mz�t^-,,�����
`�=d�`�	�I�^����`���D;R�AaS��+b����?pG����GW��G*��6r��Ӆ���H'ZA����F$�)�x�UBZDkL�"8 ����F~/|
��8:����ԒV��e��O}'^�>(�8UwJ?ܺu��^fsuPI/DI!709�%�������G������/-kI�G!�DF%��o4�Pҧs�"�8.T�J��wK*�� �8i�~�+_!���k����Ac#v���=�r�I��8�O��������3�� t���v��۪ә��w;J1��tz���>g ����8~�P�YZ�G(+fТU�:eϾug�G/������v��j�A%��J��&%��9Ϸn���w���f�up��,�C4l4��&�/<��T�%�{ICkx��2p¶"�P5��3���RG1��GoR�%l��+/�d���-��$�%C�L7ln6�*�˴L7N���Ȗ�������ƚ�.�t�\�8����������>�sV�D�M����l�?N�<��c�z���W�����_�4�TZ\繳�ڏ^J�n��[\6ݜ�+ik�ʐ�&&�k�:uc8��fN����W҃����O�{��XnQ�	�8*���D��8�B�̩����iZw�i�9^���acuie���a0����1N֓�쉓��B1U��s���=���9VGA*�	����+��Τ�;Y�1�d�`�
"ng�������?8�����.�Z�MUk�|���4s01g:��F���)(�M'��4,���i��>���]QC��Ko<�ȩn�S�+�:��gz�V��y��F�Ȯ�:����4Mt�OfhD׉�%�7=U������Z��XV���#B,�A�\i2�:P2��e*���m��ǡŽ�X�0NP'r���Eֹ�L�U��D���(]�,��9�?�*3���:w�ܽu�������C�?�\e��k�k\����3S�+���"'G�]������}J��va"Bj���+���9������.!j���\s]֪/��R�\��i�J}�Y�n����'%ʨ�"�Es7$ %� ��6ioH0�J���%ᆡI[϶W� �Md�(%^@���oh�ו\q'7�]-�T�R�pܕY�~���z�*4�- `)?�搮�R";
]��[N�-�!����+΃<:1�Y4���E:��s���� JF$�n|ss�^#��4xzJ�{z%
��S����LOy�a�9��4�'N@���#�����46p�k�n�/�z@�7�'�G
��ƖSq^!� �2���[���At}Z$��q�J�*�$\���5J� ���D�4XDJ��U�>tנ٘)H���0A�C�G:�.L2�z���H݄��#j��*F��Qo0R6�*V@��GM���ߧ�y�1�J���)�}(ᬉ����Z'��T�rm���7n_Y�o��M����L ���U�h��������B-a���c�[͎�h��a���������CE�tZNkkkJQ#�����Pu"��M���%��0t�ba|�����,K�NW�i��e���3=3eК�1:��.a�h�M��k�*��F�Q��O�B��L�+�#�'�]��@�hfϝ;�h Mʋ/��{�����R���Ҽ�u�D���<�g�*�� Bhm��A�o���T0L5J2�i��΁�
��ɲ���Yj|�HY1�Q>v��l�T�H7�l�V��*_��#}���"���&H|Ϋ����_h�4���6	6>N�(%R^,��:��`W2��md�o��\!XH��ʡ[Ʊ@���p�'������,@�T>䑎��MB�jwձc�߸q�T*>v��R��&w\��s�#0���ݻ}�6�oZ�����r	�XN>ՌII�x�ôar9L�w8��}�����wC:^�:&��	v�����_����Z�p�6���t�9�H.���0Ѣ�s������Й�O��D���.K����d4�����/^��я~t0�b�Sw}���L�F�̚���j���$�s��#�):b��cfr�yc���E��9OeB��S0f���Nx���(�o����;Y&�$|���8A&�tzN�"o����֬P��6O�E�-�X��7v[����_�����tU~�s������or7��-..8+s����:uzu��ڽ+��p7W#�6Ե��2u�6�٩y;��f��P+�b>���ي��4 �f�S���T�	lh<�3�}�����6�?���?��/�jӟ���ޚ�iqHf5��o��V�W��㠔/����A�ΰ�$1tf��8C�3ƕ�V^J��K�Y�7�ϬoS�T���q�Ox�lَ��Ob�ɕrv��,��i�=�e�C��i���������Lmfqc���/����~sg�^�T�a�ej��|�a�\��K+�)�4::��1��*A�n�={�죏>f;����2��0ӏ�q�:\�j�biZ�Ka��b�|��I����C48ڛ�S�m��Г+P�D������I����q��d�9����������F뱓��Lm�xu�����+U�´�[~wx����rV��ӕi2�$̜357}�Īz�)'>�V&��sT��g������N���\��G�N��lO�����p���Y�?��.r�v��N�r7�X�(�^4��+�98 �l �z�a:g٥���DOI~��H�G�9*�Y�:l>|y/ż���^ҁa X�*�4.�Nϴ��M����ջJ%�#�p-O4��U����mx�ޠ Et&�OQ)�P�@$
I#�������Y��(�|T+ �U*��p�lj�Y��bj4hl4���E�ZP��$��HA�A��.�3���20��{$�82L�؀��E� 9'����:�/�	�����P.��ȉ�� џ����?�D�*R��"į��>ƣT�وwëM�����ҀE�C2���w����<^fZ(�Wt����Zzk^3��4�z�1�2nKSi�*!-7[��ܡ=�R3����_
���w��ܾN���_������w����+�>��SQ�0b����+�����h�F8k}}}cck~ᘗ�r��E��������R�EN]���(:<l���K�����*p�ټHuqm;0!jC�Nps47��ԓO����D�VVN�\s�V�lL3�5b���xH��������}��͛|p�̺�iq�{fv�]'��xLt���r��2�饗��ͯ~��P{�ᇔ��(I#�YXp)I�@)q���73�%�R4���$��0!��J��O�C�	Ǝ�X���Jg�|�%dx�Y5�2Lue����"����=�;��P����G�%%��Ae��JГ�*���a�JwW��V	�_����d�I$���c�c�����n�|�D���ka��#��d���`"蜤�C+daa�W~�WVV��Ly���^���+9?[$ԡ�2�5�CU�<���|�ʕ�;�{��5��<e�0b!2�z��~�7~�\��s�0��Q�b���,c�I}����Y�=5�D7�t�����v��sǎ��誌	.n�9-��h�|��]�~��	�	i����<���9X�iWnl�������:K��\u-���`��_���C��V�;���n���{�/~:���כ0��9i�����]��;�fW��=�L��kB"n�2S˟<q�\\�~��1nT�5�d��'��4H��v=�6�G�[�p���V�k�^�(@���fyN�\N4��P�L�N1��n�'�X<}J�=��h���f.JbV����4�%����N�e��<'&[�N9��H�	��MA�,MXJ��N�N=⪭�n��qY�kW���y�3�<<r�axD�!
B��J�r۴�a�޽����k�j�����]9i�
?d;�|7_I�]9Ϊ�!� 0g�����GSq?1-us!H#�m',�J�R�0?7�8�G~��N�9�#��$��:V!_T��l�M� J�r�+����a��
���UZGdj��g>�ԧ?����1"�/<����������ŋ/��y���O?k��D�h t�N�wo�AJ�fU�P�1����|a�Ŵ��H���Aђ$7��'8���4~�eBl_��05(ۉK��G�q�;�|2��;g����0J�B3?�H��GTh�V��$��p\�i�ų���� @�"B�|~za�vl�8�B����g��CJ�>�����fLO-.��9v#��;�~o�eW�.H%J��:m[V�T�,�~�r�e�sYz$�0��Ã0��f�x"�#���ѫmlm�J9�Gۆ����}ř���4�A�z�����K"K��I+ញ���-���ӓ�T�$�j���&ס��iJuT�S��a�U�,v7�_	?
.G�%Ns���o��mZ�+(���\�R*W�]>"���IGË��Wh��w��Z�	J����˕)��1M���ʱ�����UmO�.upP����Xl2o`��S3�J-�8���ȡ�p\N�ʿa1�5�Je
	]�Fk<���rN�*�@�pk�g���m�QH�/��U�:�M;�j���3��m�LU�|�?��c��N���1C����ym�"��M���a�	��n
��8�)��%r�`�"=��2���hU�H]���h񃶩j��8H�A۔�;Di����n<�j��9�����G�UK^�-KN��}���D�:EF�4�,��۽٩N�����ȹG�w�/_x㩧�y�g{�n�\ @^�~�޽�ϟ?~�K��Jv�^avfN����yz��������4-=��GaT�U?��O�u��k��[^��V��� ;�=�|*���������?�����;�?��� �^)Vl[�i���((�K��M pV��,��{�ɥ���߽�9�T`�@Ԃ0��<y���(�C������1I����1F�����a�Ǔݪ�A��-UqT�o�G��$���Q������rypNp��g�n��9s��圜��ߪ��K�VY�<N�7�}l��T��#W
|f�Z����׿Jߤ��9�̹n��5?%� �Zǆ�.���$�!ދ���q��K���4����I��>���]]��� ����a�%H��������y"�M������:�w�U��Htk��*����H�E����_�u�}A��+[&���p�8��8����?��>����o����k�����V�2���-��Od�"�5+��'gJ+!N��M2��ƍ�7��Ju�R��5��d��|��������_�Mqh��V*���;d�i/z���i�w4��}��W��7]/��O����ۃ0��o\�z��n��0��>���g���iD�Dͧ,9la��yh�"3M�����eHuq���t[ZC�x�*��������L���l�#�FH�@��Tѐ�}^J���3.K���|{m�^�3�bs�Rk��o�Z{�����X5��s#ǄL*-���K�h�
P�\[��k{�[#��я>?�i&A�ߘ
r�*���X����B�	���lm﹥��,���Ya�@����4v��OB�}=���͍��(�����wۗ/�r:nl�.�z���~neE\`����!�t����F/,�<9�� kŊu$f��%��}���gW�>��Oy;���X�0sOgf����w��ww���v;�A5
s͉,"��oE�s�O�^��y��l�_����>�9maQO�3gf��_�W�=������>��g�|�1�-�d=}gw�ͷ����ˇ�=ZP�n���7��[���ff��N���B��e�dY|�_2�t8���	�N�*���d����R��y�N�K�ύ�,"M�n����:$��7t�Qr�3�j�}Gч�����KȜ��r�7L=��F��V�� Dk�t0�����'H'waq履U.t�lSj��p��"-�r�F��.��^��zv)O��6�;,й�j��yN�����.�Fn���n�Uf�f��J�)^�O�?�9Q{H'hR�����iw)E�R:��m�i�܃�(����RQ����_x�$�$�O���I@��&�G"K�*���8�o�B*�Z"��
��
�2;|���U�}$�mpa�@zA*^��å`	H� ��ҠK㤿B7/   @�H�u�@�dQmE?�T�{�`��U@�6iv��1q(�s�>4�%JPEà�A��hDj$(�
`D������!�M��AJ�n�SKW@cV�a�
y+������{��A�[�sx����.�i?"s$����x24�i�/T����D9��뫒���V*%�r~�.z<�qގU90�mvv��ŋ�.����t���F����{��1��F�+��x�rY��⢩���O//��ktd�������%���=C	r��a/,.���݈�����Y�Hf[�er������P����)��~���r�[���:]y�ч��pЎ��e�Yq!1���Jӱ˵�G��=3r����7��=���X �=������amF�U�V��u�qQ�@qx��D�(�@��x��Ė��"���?d_uA�������n��#N��{�Z*�'����)�2:s�H�r�C���j��.X�P)ġ!Hĝ�L��=�ͱd�"K8y�¡�c�޸���/�A��߸�t��BO��h�������"BY"��G�y���8j��pc�)�w��}�6q���4���zH9�A�48��p�о����$p��E�pd��(:T� 8 Ec��N�]�[F$���=��S8�e;(���5����P�C;������ɳg��i7�����X��6tv����k�X�R��.I���U�	��n�d��2S�����׿����/ε{C�C"a��ԹU��{�����5��i{�����Ls�_��j�5�8t�~�Τ*�v]�1B·^I�w�R�S�T'k�Ҿ[�{8���L��p+mV��q��C�n).5[H;��=�G�-�>>m&��Q`zZ/����0�T˖��S��ҫ�~�_zz�)�Ov>�9[���#��$��R�q3͂��Fd��4J�ܾy��kw�U���}�#t�Y�m��ۭ��h���$N:�A�׉l#_,��Sf~���-/VfO&Z�֊��jԺ�2�q	#i����A�6��o^�z�r��fJׯ_�ظz~��z�����=�x��y��'�K��ޠ?lt�����s��|.�&ZF�����2�T�j�J0)LMq ����>~����T�ZMb6�N��ܵ�`]�t��_���._i���,Nu+W�\[�7�#��V(���H����
}����<��s�N,�y��o9�����^��'c#-��t�i��h^�v��������ew���E�]��V����X����6����:7�`=�{���vi�ڸ!o29+t8�t|Q��,��#�$�'�����h��IB\��e,;�d�����m���@�Jqu5#~�����{A�kq�T����#Ц�+��������a�#�s2ri�X��>��0���FL��շ/]��zj�#������b�p�����I��HX�d���>N~ED��
ƾ�7�A��v��ۄB0�Ț����8q�F��*��7�@?����=6`�^���3�M�u�'�@d� ��	��Z�R�g�ODL�s������FC<(����%�^ �'�Fύ�-TZ>]GaK�qɄbDEH � 5��A����z:J�'0$��d\J2J�3��^R��y�QI����,2�ۨT���!`�0"��-&��G���ACz�O� �@�(u���$�s
/��۹J4�r�?�Q嬳p�:5U��!*��/�f:�c��ŕ����W{�����j�ԭf��i��ޣ�=����oS]2h�󋞗/+�mI�/�s��c�h�05bM�R������7��a�o�:�{��#�ҏ'�QV �DWz�*��'�㚅"}=����Q9y��+������
��@�S��s������Z�fujjy�Y���}�
'4�P �B��V`]�lmnn�X�o��*�ڐ)}�lb��ȥ	zI!~�����tn$1"��J��N�k+�� g&pI#�&��z	4p��|i4�ӑ�/ˏK� N@��GG��� Yv�J��u�����_�)�K ��N�HXEe =����$w�TO 1d���fى�H��w �ZK��q�=���S�zGN��|7c�3�1%(�9��lmm!�.����l4�5�ϒ牚I�>=LtV���.)�Fj\��hDK����o3�7��}©�V�?${��R�t �	 �<y��q<��9�lj��:�'�f"t|u�#u�!�����۷���t:����˗߾z���H�q!���!�9�HJ9F�Vw��lq|��m�\z����ˮ]��;L�Ӥ�z��{����}�h��f�R�p'O���ڧ3���mٔ%�C�G!'�K<HY����X"�
�4�*\o�9<h��5[�A�-�����b4��(g�;Teo���2*���X�Cv�h�0J}�NA#��=�8�8��s�bn�d?v�dezag�S��F$g�Tv�����A;lo�>!�$�0]%d��9�N+o�+3E/�أ���������ܬ��~@w�ƾ���ٱ鱸�t�|~���ŗ���C�m��0`�o�;��h�v�����k{�wu-��*�KD`�NNw���GODC;
G�e����� ���5��\����3U�����\�F[�e���1�#N-ct���;{���D��q]����y(�'3�^���4��0=U�v��o��z�$Y��o]�˿���Ζ�t�2Fwvv/]zs��I�+7�ݭ�Z��^��䫕��/��/�E���n2�@r��9������?�������~{q��l�X�6�4�i�N�ѭ^���Z��Q(Mu�݋/��/����I7�)tj\�.G�#��J�j<)�S�;�11xQ�K�L�ǩW:M��ɇ��ڢ"�AWe�,��\ײU�^%_��f8n�3�x@K�������ͥ�y�x'fp;6z^�j�Z+�f<�K���4F��A���+��v�x���<QQ�LT��f���z�+g��)3�&��.7��hJ���4��
�芃��Ѩ���P�N��K�U��^��؟H�9ש���PZ�%`�#Xa��PP[F!;c#������0���]3�5����%b�@�jm������ ���s�m��������)4��?�oR$t�G�_5�i���x�n�=����Rix�ɨӾ@�xQ3�m�J��q��Q�ą9�����lWD� 4�D�hqquV��*�y����I{P��@A��&|���AE�5�T�2ITP�+�'��������Y�t*�5�(}�\��@D�5*r�8
��,�T
|	�±,R �Gxw'T|L��h{{�v(��>�eR���R�
�]onj�ˍ���s>s�0Z:��%��Q���i��������������i�	����Z��/���ڻ�c9R%�GW��l����
^!�/����*���?2�Bzz|�� C߈4W�Z*̢r���E���9�[�Σ`��s�jK��.e{�7�G:���[,ͧk#�Ϝg�FL��r��L�D�MJ�ߧ^�
���<�w �w�ILU E*�=
�|�rg�D¤t�_��"�<�x'h��
X~%��?V�eU�>����-�h%���`E�9�������j5�,����_h-9jq2v�5ٰؿ�j���Tqw�'��eFI!<HRB��� '*H��b?�h�B��-�8\?0
t��r�7M�!��0Ap!��/I����,:Zx;@��H�k�M�Q�j�1)L��#"!M�g��PM��F��܏V�Ja.~���"� 0U-��?
!���1��T[T��4����Z��FQ�z�V������޼�v�Xtt��\���Pf�}��[]9A 8�G^�pokw�i9������v� �3�8��:j5�*��6��mz�J�z� ��%~K����g��O�Y]�^����.6q�Ly�,/����*�f�1��j��j�F�ju���i4�'WWW������I���^ȉfܩ4V�����	��2lBW�A�U?<�P�����_����(�n�~�;�wr�ŕ(1�v�����П�?��^�S�Z���+6���.���'p��ŋ�����3���,�V�H6�%*�K�؝�-iDr����k�g�8���^�3�SCOL�<Ik���흽;�{[A2l����nk�nm-��ӵ��奇~��g?���ۍ���h�:�\ը�Ť���o~k�6575����Ko��l5���H�-,�b9;�������?�����Sg#zX(W��A޳�x�z��s�t�C#�X���J�$��'_���v�ν��z�ҥ��0�Bn>�E�P�~��o����7Z��ԛo\���}�����_���n���>{�R�4Uay'�L���5�_��ҏ^y������yg���o}���#�K7�_���vsn.�� M�6�×_~�w�wuӹ~���7����I���W��X�{y�~�����Bv[79�@�n�^�\�{SV�,y��y{I��R�+�~��܎X��K���]����h�*�B�C);@8�6�E�ghrF!�#y3�#=�eʙ&��a������N�v���G����-y���N3hCzvd�[�������?�c���gWO�ԭ���������Lc0d���F�~��� ɋ�9��]�حN��,.|?0��VMB��(��J!& 	K('	8�򊽑���`Q�����W��j��z8�r�����@@��t�6V8��0.�Ҵ��W9ܜ�KW�]M��@�T��[���Z����	��A{g3����O�{�kঅ��>t��8�=gcH��`�ߓ�=�F�ѻ�-�
t�'����K���1�B:� $\��dz�]
-q}��#��@8���+�#���D�OJ��n Hahm�@Ʀ�c�� .IQ�C�z��C�^
|!z�7ҋi����ᡗ��SSH����T��^�[.�TO�է����65��Qo5=/���j�5F�#�*l�b���ǵ��L#��C�J���\ͨ7���k�ȭU.E�H3��g�]�v�_�ۡ����>r��
-�N�5�����N�hp��
�=Z��X�~���G��V��D���4��O��W��w��r����^y�B^�����i;ޠ��6�K�T��e��2sżc�Q8�;US}���D�P*�lB�@��r_߱B��j��[�=��J��aS����+������7+J�x;G�m9�vQ�3n]@�R%J��HÑv4ȡ�٧5W!=���k9Wu�����y�+��V/}���(66�בtw��m��X�tp����qv���d ys��kୠ'��OB�u�qz��Ӄ��Ig0*D=R*4����@*� � x��$�D$�5]r�,�A �'���k��7�4�Q���{\A�D�L�h�ANE�Kg�}=k����p�D����fjt�01��aCF�n����իW��K���W����qJ۠'�����Q�kЏ ��k�]%�%��Y�l�l�Pjyʲ��v7��>�����a��f�rG&sŎt�[,����mn�C|���a����03��\GB���o����YI�<�` �M�8�>Q@.�5�Q�NrD���N��c�=��G�����W�=�wʝ�~c�`inv�Vmk�!�s@���ۄ�	��@�])j�E�0��Q�é�B���QT�ռ�����;�[��v:N:�rl~v��X��أ(͛�T�j�N�Ti5���fw9����wZ^u�h�0�͑A�+�C�����F�U���;���_������g�kɀpA�v���W�^���~{�݊CLto��qXGѷ��Z��J0i��-��d��V������o�����h�l��MLc|�N�`�$L## fM�Hc-f��������>5;����3�q��z+�탳�~��o|�����ʮ3�;�:{��4�F������/��+�&�	�Y�\z��+���W�i:Z�u�*6?R��(LiHid���W���_�.�<z�*�0�H��752(4��� vUK9Y)V�1Ȇ������J��A�#v����l*6�rt�B'
�4\hQ0y_��2�j�(M�C�e���AH�bA��s7f�M��[��w�8��%oz����v�ڵ{��F#�H(�2�0���Q����g?��g��y�G���������*SQw䇃(j��*aGh�qi#�m/M+�/���z��������p�����rp�.�s��=��Mr���x n���E$���1�4"> �� p���$mgM˃�E2�������Eox��B�D�Vj��/�BCE/� �{�Q";��~�:������u_t^�%���FC'A�0�$_����BQ
��
���z�,8�=W�p�� \�M��1��'K��<��R�I�� x0�'�5��a�K�!&Z����ަ_��͡6Z4��˧!�<E5��@� ����S�Z7yP���F$�$�$)7�C�n�suV� ~��#�6�]ǆ'^)����&���c��+�w{��y�6�ILO�aV��/܅��L����d�f������믿����O~��ӱ�K�1��eY���i�9s�����.0s'Ҕ���Md�p�S�WAv����}��Z�yX�;]^^�g�������?����~��29.����~���8;=�rS�a���^C�/|
�>8-�$l6����ٳg�5DB�����8�z�Ϗ�V�NǙ�x�a���I���C���g�{Y$ل(Ԅ $mt,3(��:��tYŋ�Yy7|?q�]aww��RR��A`�VHN �eD�Q��g���H��yс@�G��>�%8~��3��C�����ټ�w�L8�t�!�
G
�t���w��T)·��s��80QE��D��Ȗ�	]eUh7<��Eg�[Ƚ�	oM�|�xV�O�K�=�B�;z��8��{q<y7��}p%���lл>:���P�/,,���%���� -`i�r�E~y��`�!������I��Q����Z�׹E��j�,�)�DKY�GU'zӼ;w6/\x]���b�Z-�[����JmV9+�9Ê�X	��N� Ɵ���_Syd,'�ou57�������N�u���|칏�8��L��Y|_������ �9M��M۝��G��Aw���-2�H��o�(ҳ郰g�4�͟j�kk�b5J���Ny�l{^0޼}��믮��J|sy~N�j��b�9S�Zo��)�j����o��[�˗߾�㿹�8�=r~�8�������4���R=��OWT�e	��pb�vG����H�>	��q��l���N�ܣ�B�c� W�'�s/`L��2$���]v�&�dT����3�hLA<ր��d�&-�T�XM�̒��ՅL�t�\���%��Gh���#S:?��@�oǉ���P$'��?������<eb���{�X���к��o�o�h~ֵ�\���h��֯KB�����m:F�]������>���9�D?{���ˋL��S"�P`�R�)`�GF4B���v��s�:w�a�JFuA��
v�uF�HFTz�� �Y[!B�T��x�y�z��Ir����X�.nK1Q"� ÖS[� �G�o���˶���I��	@� kk�S�	n�lP���v�F�~�)x>h1I �#<d�C@k�k�W -�*&a%|��EEV�(`xB��ؑ1���	!�� `V��H�.9�J%7��"{PT�pM��P� e@@v��`���	_�̝^I?ӻPpn)QG�
<C<�+"�	�
8�/�\�� �����&���e�ױc�N�>],x�<�ڌ����I\Q3sfS�뵿��<=������_�Y^=^*M�.����EZ߃���n�.�Ga�m�o߾y��%��CR�'�����ꩺ UF�%����� '�o�=AV%yr\+sO��e���[/��"�,z}Z~t�Ã�n�?{��G�{�,=�F��o~�������*��f�](�n�]��ǳD}�D@� �M]���Ӵ�nܸ!���GN|�ZZ����	�t۝nw��/�s���"N,]4���aS �*�X��Wt��T+I��(����}J�� ���
6&�8"	�88�سi�X��i�s�޽{R[�;�r�ɡ$}Z0f�����!+u���F��waG��$JwRy�^���N��;���DH<�Y��#���>�|6f%�<~��[v���b;����!f��!g��Ѯ��ƻ,��j��m������(�M�R����R�l)lv����]N�T�r��Ѡ,���bB�Q��$4@��!���$qښxY'zbc��we��;�Vy�GA.��6J���Y�U��w;C"�[tRr�-Ѻt\qֽm�vQa[�9J¬gG)u�D{W��#�:�����n�[?l�z�A}���{��cg��,z��mF��U���Ӊ����R�^�z�3��n�߬��B�νd��4]��2dI֦J�s�Պ��w���7.�?�����V�oݾ��Gy����`�5:@S=7��)M��
��{��[Q��|�«^��O�LM�@6Q�e�t�+�^�;�ߝ�I� C���a�+!9it7�����H��$=^���/�L��^E���������.�c	O��'�F��L7��[��If̆�[)�s&��5&{ژ>q]\�2�mb�cd%C�?P"$���
:��r�t:d��5�vh���G���i���U8��agr�# ���o�M�]��b��Ff�~��?C��Z�*!5�YZ��B-�kw6��!К'
�S�r,n����7������J�b�����=��SO=�}�*m��Zyff�>�w���6ݲ��B�UH��@@�-��2B|D��K���!�x��X�8a��jV#5Bp9d3�:_*[�i��=�C�"��+f��Y�2F�Ξ���y�8qB���ᓀ?,�B�4pYd!5����dR�MG�6��p;����Ǫ'���h�'4\psJ#�<� F%�� z-���K(��`P��� ������}�x��.�&0At� 1Y����Z�FH��%�f	
�3�}ѓ�,��g�n~�pTw2��K*�q���bT��c���:����4�;�n��h�D�zJ8nqi����%�:�fol�3u�kM� ^1?[�v���޼�ȹ��j�A0H"a�W�KdY'O�^|�����\k�%�l��m�:}�~�I��~Gݦ��G:)�L��$JYSQ�%%@��00���l���~�}073M����K���t�?�+����8��-b?���}S��t��,e�SV�B�M@-�Rnoo߽{�ӟ�4m%����b��x�٦j%�Z>y�����u���=O��`OI���"�$c�y��F���į<��0a�ȘE�Iu��a�H��ą�}���ׯ�J�G�O��-�w_ߣ�
��&	Dg�&H�*�0N�qB��<��v�]�-)�!�y�� 9f�ȴ��#��>�C��r��D(7�N�&8���$}�!=�z���T�=�r�Bg%k��~�/����dⲹvع��)��37B[����~��li΋���%�?�Ў��h�p�oڋ�]%Ԥ��*O�6�e굙9�Ԑ}��,'��q?���n�|�h�sM�pZ�7�MUKK˳􊛷�[�mGA��?v��z�\������-�4�A�����`p�ν���߿�޺���&#���Μ\����;=� a��"�X��Q�Z۝N��/LW�t��,���şE�ޥ
�H]2	�B^(���������������y����F�����>���rz�W��#�����PQ���^F��na��˪6��&�&M��HA��33��zd
��wN��\q1F"��d#�G���)��S��ji%���#d��Y���Y���<deqRK��5�-��o(�dUh�L����]�b]YRCO��*�W�z}$;W(���(���F蝞�4���q�����q0  +=�)I��9Ģ�|����8��S��zj����U��˧v1��C�����6C��IBM���;\�bpӞĤ����YFlv������ȣ`0�aG��ų���ԳOsAK.�G���ܩS�J���`I#����R�T-sV�d߯��j�t.J�	�N���)����	��[�o��ƈV�X�.U��;������8�I�l�x�F]�DaC�F�?J\�hA@
�
	*�d�d��k��&�9�+�@�P8�"D�C/&�F���ڢ��d�� :b>��P��Vd������Lz��јQi ����W_�!\)q$<v�P������o o�xt�!h>��b&nl�Su2h�#�
�p&J�,G�� ���������p�H�a��Pz��)B`�>�g���A���]�����e�8A4z=��p�F*��v�M^�:��ک1��K�-��^����ԧ^x���[7o�9}q������h4:����R��8�T���[o�q���'W�2=��Eۿfx�֭��Hl1ڮV�Y�4Iڭ�l[��Г�R�{b;�����#�j͐�oܸEˏF��lN���(�üe�HTw`���~zzJɤVJ8��(�%�Ί�/�4���3�'H��%��}��I42R�;�
�B�Q�FS)"%�w�l";�B��H����M�'��7oޤ�gϞ%J�_��&ݍ�3B�*
��s��{����XHB�E����Hr�����xW6؂9E�-n\V�J�
�c�55C�U�ͫ��?z��f���=�N	��T�{�>�;YD6,�@_�Γ,%)�������zѻ!ݱ�ЃJY��[�!��_9n£�	��@%��2�����m_�d��?ː7E�;���w�;����bG�x%J��nl&K]+x��	X��b�25�������0���߄��v���	�p�h����9�%��̜��s��j��w��N���o|��X�̛���N�ӕb��~/�f��67_4�E�8U�n��a��1��c�z+��e�������D}��~�d�\ۥ�G��kw[ͮG���]]�r���a���/X���M��x���i�TS�b�1�3L�9F����\�R���G>��k�R����"�C;���_�xZ�OR���}��I�,���d��G�NI�W�X�詡�
��H74K�E��0	�������JGYp����x�(�5���y($Q9��A�#��p^L��?P"4>a��Q�T����H!���'��6ɦjI���CLM��%�64Is�镏��3_�׾��/85-8�/:��i6�~��Q2j�t.�>���P��w=$�],M}��~���c�?$��`�\�FFA����䀹�Y�^�88�:3pyw؍�y¸A��a9��`��hC:� ��@w��p@
���#5<�����̍ ���"���5(G�ɺ�G˶A���8���ʨc�"����OH��,�����B�BOt�֨�G*^)���jI(B93�v���t���.R&P�FC�zO9��qYȸ���*�R�2G�0^L=�v��sZr?0��C�)FΆ*�4!��;�=�����$}W�^�m=;,BTP��qA�PI�A��xPtM6����	�xj��4�^W5!4�􂅅Ֆw��'"9ݝH�+��4l�� VVV��#W�w��v�(�TKe�1o䞭ʱj��o�q����k��e�6�%���������;����s�Y=q�V�[7��֙ӏ��~���](��d�V�T��W�� 
��k0`1�G9_�������{[��2�v-��]f���
h /���肥R��f��	.Ьiz0;7G�t�}0�G&�$�P,j���0J����\نEr�әCG���.�ݻw!$|AK\����O?���G�N���Ů��8L*;(г�U�'M��4�=��}��	��I%R ��;��25AGs��E�ܹ��G	�:���N	�K0$�#\�m�Y 5rȪ�*��> {q`ey���р�$rq����k'����9�������f��dה�+�n˲�#QJ�O�D�@`����VFl�H1�n ��l	�D_��Iһ�ShX)�[�C4:�2�f9�Q�`��8������AH�a��ͺ�i6�4%����M��N�xR��*����z0Y���DO�Z.w��0HݜCf���ݺ}��E�J��)	.w���ޅ�c+'{����[d�a�r�JY�����1�<{0�llmz�h��ٹ�N��`���Փtxz�Bw`��+B"	m�D�/�+�����
DP�"T�c�RA�}��ǏECvH̢�ř�Ze��K!"���x��s��n���W��;�����\1G��К���t�eƄ���a'�[�����Ѿ���w�cZ��.��k�{�q�%�d��cB�._WRQ:&3�&ҼP�I��K}���`1d�I\:j�ʠ��J�qFd����զ��&�%U�:��B�(�l:Ex8���U�,�4�w�4������I+,�l�45�H�7�J�D7�Q^IS"��wv��o����M��2J�Yv�Z��Iε����/O�~����R*�!D#����5�K��p =ҹ��j�6h�Dd���4�VV=7z��+�,Z	y7Of�'���̎����C � 9�dk���D��E)�$7��㬗
"@ѿ�e����2i|.�`�5Ŋ�J�����
� �H��A�i�����rHՄ�����+���D�IJ�#x�eA�`hE�	 �ZQ5���H�6�\
дO���+	��Y�@�m���� �P$�� �!eQv1HV��.[�0�*��C�����D��0<��Bz��`e�͕�VAb-�#�B�����"ޠ�t$�MMM	A6#H�#���w8�1 ���r��6&�x%=��W@��������)J�Z��e���&[#�]*�\~�v���g��.�lw[�b��zl�r\2�:��0;�6}�'>���}����4��^;Vs��{�6}��u�X��f����p�~P��Q�"��45-hr�l�����$�iu�}Pow��I��p6f���E��� 2L��M��)D�$E[�u�����ؠ١�Bj	������&�8p�W���Ve�G�����J�l�4N�������P���r���0�4���F�%��4�B��Hu��đ�=����HEE��J&y��0������#����_oAY���J�%�)���2�\%��%��z��Α��!��U<{�O|R$��ٷ�OD"[O�M}��?2�,� ~�<�HK�lV����W�V�j��j;!qr!`��bN�'�Mp ��E*�=�
3������,*���M��w�fS7�G���Ry�(Baq���[�����Q���p���m�)Q���`ie��?U.M_x��ntn<��N��Չ�7T��4�
^�Tԍ�;��Q�b����.�s���f!=T+��~>
�e��-�9LKwrt������y׵s�.'�G�c�xq��0����1����]NZ�ix&��C߶��R�*/�hP�V�UN�o6��V;��n����7m3�=��T
S����p8aS�@|�(S�lfZV�"��1�d�2-�]�u�H�ٸ����E���Tɐ	���kԪ6&W�M%���.3%�ޤx2�F�<��sN��fU�D�����Y�/�P.�D���G�`�uē�N��(;�1J:���|�Y����Y�	��i��� �!�����h'���m���a�8��s��n�N��o�����hdXn����|=�5�aۈ���Y�~/(rC�ۥRx����g5F�ˠ��~�`�J�PU�<��ٙ*�&AN!�]v*�|!+ &&9��IR���`l9]P$ಝΥvfI��K��2h���M�#Tzzf����憘�v�+�)�G0aL|�]K���@HxJ\��6�oP~��gx���Po$�MhR�C�,����T8��իe�o �����>�PB�沣""��%zD"�%1@�� ��4d�R,$��t ��:�}��W�fii	�?�pB>���zf��������q��K��4;;K�:88�7��N��S���zf"7�������f�9�l��'�Ԕ�5BƄ���� 2@Ϳ�0�CDt-y�����֕�����={fin���v�Y0���ʷ���w�֟|������W��/^��w?���F%��r�NA�>�������j�=�l�M�+�n��61s54�$"D���z��1ŗ-ӥ��8��{óg��9<��3333�es�;:C��3����ǎ=��V>7�D�nܸ���������/�z�X���B��ē�i�X�4S�����O��Io��ܼ}�6-���Ìg��� �RB`�D��"O$&����P��z�+K�.�@�O���Ò����/b�<^�8V��fpm���f
3��"b�"�T:�H7$3}4�����YɁ#rgؒ����%s蕴*p8��=H��!�G�f�'��������wE�Ry(��C�w�QG�~��ȼd+�|f��{i	��8�}5b<�a,)pRY��ZV��]�����k�K����W�p�Bj
�����OO���!р�p���#��;݌�9t�EV��Au��Y��K�N=��Jm��J����������ܳ�<����Ko�y���{!�/G�P!+��`����ҨT�y�&�08ݧ���9����|�<3����WZ���˹^^+��+[�V��3u\[a�$��Df��`t[�n�I4�G�u����.��X�Z3L�Ь@5�����K���/�����p{s��S�|aR��+�-�2F���'ny|�� �����әr����J�t���	�U�GE1tM�o�]x(�']�H�
R��8=)�ǭA�����Hs�&u����W�,�);G`i���K�H�p'���"�K�Q�Ed�3X�� �a 칬�:c��r�?u"�G#���k���:����4�1S+��Nd���� ��p"�;�2�!-��P�{A��t9�I��C˃tn���(��$j��z��������?)�3QJ�) �M��v�fR��L���x��a�-W��if�b⸆?�٫�_��W��ի�i�?j5[{�a=я���]��a@D�0GA�V�u��h:-�\�*Ŀ���*K�bTPH~�h1g��#�I�s�
�fT��Й�;:�/��=�gP�Tq@{DvI�y��(ͤ��HԺ�����.�[�h#_%+6L:!� D/G�x	j�P/���1S�>�E��h��Z�50�x�x�:y�$!0T��z�*䤡6��x,�swww~~��JD��$u8(1#o��U�DK�!Qi�)�c�z����a�91�����C�&\� `�Y4�4T���E0AhCD��h(c�x Q�����["��ݨB�D=:]H$��NL�3���"�@H\+�Z���90,8����k7�͙�g�|!Nt�+٦;��F?_���[֌׸�����*x15]��nd�[��k7Ϝ:SI���Z�����@����U�3+����ۿ����2�H�Ce!��7�&����
�R�-�� �4�-��ʩ�K�j7ϟ;���:��;��c��h֔._B,~j�Doz��������q�M=vb#�@hnmmq�yn���G�_"?s{{�(��N�8��SO�0�?�]����F�?���O?�43x�@��!wN_4$��L
6��B$1P�Kg�e��|)0s�#LӼGd3�{��t�Ŧ>��vh�T�-%Eg!��	SK���0��|:�{LG�YC�X)ņ��O��4�9�ݵ�|jZ���d@�u��GZ�Jz� �Z�#�JͤOF�ܬr��6�.����D�]�%=d�lib�#G&�Nd�Dӄ"�Y����B'�H�ŀ�Y�r8W��H�>�lػ�Q���`�.S9������ۡ�uZI��l1R&J�0��G��6SGsR�.b�������.rY��]���ix��💐�ޯ!�@�Y�3)��&1��_����mee�����"���3t&a�
�q�}�2˙|���b��lt��-U�l�ιdi�0;�Nc���Qj�!�w�U#u8����V����,w��">;㐎���y���入�%Cw|�򫯾��6+Ӑ��Nh&&��Xnj�p]�p�a��ȶ�,��#��ң(��/~�O��w�쥯����v��ÿY��fW��.(�g���x�t�����6����A�}�杫7��u�g;���I���G��&���j��lܡ[(;����s�,ff��R�ʕ�t�z����>�Bu�k�ǵ�R��l}�!-P��ʅ��-{��6��fyq���4������+�q8R�[}OU�P�e�!�*�<;�aſL���HXP�r�����~Vd�Z�/ǿGu����XN)��Z�_�����/���ʹ ��pU�r� T����SG��:�Pk��0о�O�P �],�&n��n�ZH�i�4�-:5YA�H��׮������|��շ�̘�����'SA�Ԃ��[J�$�{�����9�?4�M�$:��K���x��Q�y��������^{��3�]�7�ѳz��S�N���ַ:����v�}��0
�U�6����w���{���V�pΫ/T�+Vc�զ��=U��$��D. / �e����q����^���t�$���P2JA����4����v��zir�+H�'�;��� ���8)�m��le3�O̌�&E� s`h�*)�����y��pGԟ܀��1ږ2�БL씏��?�8�&�L?h�/{o�$�}���=����z߻��  � R��#q�k8#��A{�?�qfb"Ʀ��H�$�bH�)��IA �F�]�վ�v�������� ��d 
�U�w���;�w�c&���ϛ΍��>�����E~��9�[��ցk�="��!'kkk���y����fK^)=�
wG}������N3�9Q��8>�[�5��α���ŀSӴ�k��l)�r F�3.}ۘ离�p�!�I)�TP�S����2ce�3;5�}G���2*��{�ȝE�G�)���ͣQn�w��^o�ҥ�q��o��5X�\|���Xk�m��6~��]��#vdЂ����A�n��j���@h����8�viqo�=�����$U�	Q���^8����d\.�J#�Q���v�<y�d�[������+{J�P&�+C1�*W�Oeey�%CRJŅM�)�1KC�����E�$:��qv�3&$1Ő�xQEN��C���E�����P�<J���4/5 �cd���
�S�䕐�K��n+�*���$�W���'����'��9e^��I�A,Q�Z�����G�%�a�,��Iˑ���]B^�^c���a,���!
��Tݣ0�0���'ZF&1y�u��9a��8���S*U�n���Gǁţ�Nז�⨕�P��c�!a�?��OA5A!�^l���!�SSS�	�a��#-��©ԥ�(M)AV�V:�<���A"��W��%ݹsJull�UJ�/	:wA�իW�o,\�<������x�iB@l ���a��[���z�*f�i��`���"ObI�~����s�x�Z��NՑ��Zd���J�Q�6=_�ת���ݢj��������q֏�p�fǅR��tL���l�YX�Cf�L"�s��\;�us��ϯN�7זV5����;�7&�OV'g�,.�ЙC�}�$�Y.<W�뽅���~������<�I��2q����x�/5��L�#N�Bq:e��Q=���cy�q�Ń'O���_~��LFN�����^;|���\6q���;%)���������������۽���|~<�Ю��{l��ADmY>$�8���8�P��zQ�sh��AA��Sɳ<1�P����o�O���t��;p�^X�+W/������vd�3m�G���g)F�l�*�G|^������?utp?�NV1�2��`P�3�J���e|�S��iBN�#�`t��-�^#\�}����A�3��t7��͛7�ٔ�)*_�c�J���]�zr��c�0W�0�����'��S�x���?`ue�I�kD��U�Ņ�c�wE\�j�cYfa����_�\�Ӆ�Ѳ5K:�1`Enܸq��	����-�E`�F�[�u-�(���.��Q�Q�{��!,��3v�Ӎ �N1�Z�c�I��tG�L��;K��a����?�u�Q&�5b�g�I/�f�H�>F�D�1zgh
{�&RՉ%��쟑 ���~��h���q�C"�IZLY٤[/������;���s��?�g�@#�u�O�-6�֠���4M����AkG�!�I3OhK�2@ �u��5��"̳(M�8a��i���]��{����mlo��օ�y�Vl�U�eԀ�hCF�,�j�����\�å�w�W��s0.�N�S?Pf�b8��K.{�8���e�u$�8��V��la����W
�	����F��:�X}JӐfU���h�QԤoenI��i�&���p�L"�����F\ Q�NX�{g`�tdZ�VjZ"Nu~1�8��
9���
e�!�zX��k��.��+R�?
�0�P��M��\VF}#�N2%�F)\Xr��Q�%K�\(*a��ݩ��>�振S�k�[���:��}^����0⻏P*���گ]>�O9��رc���y��5r�X#�HV�J,&��SI3�XV.QdN�k"�"�vYb/���g��ʊD�#Q:���P�Q僚�+���Tkvu��q}k47K��~��y~i$�Z��tJZ�[�?��?��o�rw!����S���ԯ^��-� >�9�'\vv��N,Վʶ5�go�"��ͭu��lQ��o,�������sM��
�]������O�z��s�3��M�\-޹9p����J�����Պc;�qRk�۳�[Kף��~r��w?}z��?�F�B�M��t�^��a�~H�!Z+�e�	kw���ȪA5�;�c!`*a�E�^���ge6)TP��z�Z��<�!�����v�8�$�1֬֬���p���m7��H�Tz ǩ!䇅k�b�l0�uW��L��c��{���8H͡�3Q!�"N�4�ee϶h��6��`"PL��[�X߄(��g?{���ڶ���$�=����fʋ��uMv3��±1�@����enϬ�z���-b������2AҶ[�v�,�m@�@!�}B�@D_P�i`�j�w��p����ױ�J�@��<�:IL�=��s�0(qeԥy�>c5���(Q��Ng\�@��i�b�"l��ܜ���"�tT���
��T��ٕ��۷oèb7�5����T��ߢ&3�$cP{��|��h�߰\�e^6�\|7~��)>&^ '��3���u��R3����d��44���D!�ð�,�a���g�go��U0���pm����;��^Ib	>8}���gUt%+Q�hi5�a�	}z9���SA�q�� =�[]]���1�l��)=]�_:�8&��1.#����f����S��V�W�$~��o�ɟ~���K�k�8���z��a���������{�L�=� +���WJM��bF�Cy:��a�K�Iaږ|�f��~��ͭ���ȵ焁�o��|�w�wI�����xFG�Ž�研���ҋ/���{�.~����/��/a�yz��'���-D;8��/B��3����k����Ei�kdg9�����z��U��a�n��w�wp�A��d?�G�ڍշ9KT�ΘI��.C�t� �i�8ИጊB�?� ���8���~�E#��J�)�ɔ��X���&y3K�+%�5\�(�ݲ`��� ���a~��i)�ܰ��Ek4�Fh<L��U�]Q��>0��+�m��`�� dq�q㆒���Ż.���.p/�����Z�@0σ�d�J��m��Mb*p�a��q�p���"+*$j˙�IL�`����k�UG5@Li]�r��]��i��wS�~���[��>��iZ�8m)j�~��Gߗ�Z�ӄ�ݼy�ց����X3/�0#T���L�N}O�X2k�@�R�fL��W�5n���p��E������x�U��V�&�S�|�V���@�#����A��ڞ����@��(g�P�<���4X8�z�׍l��_�=�s�ت~3���3c���.�,�I�Ij���q-'q��N<������&�'[��g5�A��zi\8)BSP���d�I�#�|��P�u^-�.�K���-�N��D�ǐ��,�z���{o��&Bcac�C��W�רyF�.�d@�����j�V��F��֨㽰�a�����s�����б#��lmu��h5'�V�����\~^h�}ѽ��U6*�G���3�^�i+B��jԽe
�p�Ӿi���pl�K3��/r��mL5��R���T��reeiT��1�<cy�b;>1v��	��f��m���Ȇ5�2S������f�� ��K�Ns����Mţ��(��{�W���!��C)�迖��B��͂�I��%�)p��E��#�
�Bɹ��'m�c2��X�W\*�*�δןѣ�cUf|�\f7�%��Xj�����^�cћрJs$t͕?��P������$�0���A�1
a�[�#Ëō��[� j��F�M�O�1�O�@�Ņn�TD\4\�2C�d�(J��8��,:�T�����	-�p�̙3��x%��U�c}�R%�������35�
�Rv�ӄ�/Mʜ#5��i_�|����135&��~TdN�%�P�f����3c���c�z����c���G&W�R��ʄ��]��"-�#�8���c=ǧ�*uV�k_��7��M�部�-3��^��SO=��!8�֭[���w��P�O�F �o���;ׯ_�)��t��b��%��dY��\7��Xg�"3x����V�����5%�0���|C�S��[L���-,���B�q�Hxa���I��p�4D��z�IU���w�sR�I�@�+��}�v5J&�!�Ra�5w�y�2��>"�Z�S��@HY[X�-ߩvCY�|IUƓ~L=I�Ö#�r|y���&�>00P�&�q��	���˦@�����_�>��b��b֮{��+4!������\k�\42�(Y?l�B˨��mE�bvK����Nj5�T.�|4��ÖN�
����*K-�#�F|���3��"�U�L���ȑ#DB����L�R����;c�Ӣ s~j��X?�+��x�[�yL(|�LZ��Z��2(m�b�S�+L���;�77�I��DAƱv�,�H,VX��oL�LD�$Cª�ꇩ�9�ܵ�?����왜�l��( �i��5��	�$~�ޝ�3��I�Bh�Jnf% ��-�MҬ�f�gwI<�B����D�aU݉V��<��An|'1D*pZ5����Uk�f��_��u�d���V�aVj*�]�ϡ�///���#���
g�&�4�,�=��I[ZZ�ַ����~;��+X�{A�g�ʤ�\*t���y��s�x�p�
V�V��'�83����|�?F�����Cܺ�����	ư�[�^�B�^f��e�r�q�+Y7����Lsm�W�5|V�r��Jlsl�J�|�ϛk�7O�t��m�p�B��sr�Bwt&���V�IC"1Q�Y��=�jIq�����gff�j�GZz��,/#����`ا� J���U�LY�*װo�>_Ǯ�O��R6ѐ�ED>=K=���3"�3O���*���9WX3O�sB�g%��B�Ӫ�r5u�2YE�Aѻ�� J�d|���Q��l����x�[|��_t��bHOr@*�ڟtxF'N�ؿ���.03}ĩ�ViڒR�+��s����ܜv^1����6�"��������2a/�x�δ��B���^`�b+ă��Ƴ��,0� qit��"�{?Fs��Ý��`y��q�ܰǉCr9Y�u�֨bm�D4�`��Ym�j6���>r�΁f���KU{�����W�W6WV6���H�
�x��=�:׫T�Q��y�۹:dx�h� �陹v2G�P�8�ヱ /ͨ��WUV��0!��Mn�h�%2@���ƍta�8�.�+n�7�|��W_U?��Hv�	�:*�{�a�7Y��e��r�26�͛7/^�8����I_�w����D��� ����h�޵�!��ƭe:ګ,�Z��d��L�e$1ǁӟf6������Kvm+�7�+�k��8�N��Ũ�*��l��88�S"x��s`1�)M����HΜ��s�h�{�[��[ը��O��>0׹�D���ü�޽-e�F���#����}�\�5�q"t��O�5᭭��a�9V���l+mB�Y�����̼���^y�._LmPA1�B[���垟]B���p�ʕ�rB��)]�YL�3kS���Bi�:ap�]��d�yjf-(q���5��\�����}qs�9�L���;�J]�2z��|�� fXԶ�LJ����v���MB��IcE&�	'�Zg����8>�';B��	�C��*�J���8��;���\OR��t�f(-��a<.:EP �ocs`RPy��rL{л}�������	�}�h���fs<ꈼ���Ն]k���%�wa?��^!�"��o�ϭ���QC��"��Yp��<4�n�	�t��,� ��p]�b���_r��Ǒh1��`Co�<yr�޽��
���f��He��j&��my�|��-W|Zؙ�=f^yltE
k�6[�Z�-��2<1�ibJ�i{޽�*(<?i�|��G�!�4�p��u�k+�k��1��v4��s�Z��!j�]u7B���S��EX8]��p��ip�=H/�v����*��EC�2ٹVn�~@�/s��:C���QR�*G�eT��I�i�{ظ�����i��y�Os{�n�u��x�z75y�����Ҫ���T����I6���xb���Gs�:?J��lie���Ƀj�H�@�^&/�I��u�.0�С���"�L�'���VRl����ѧaW	^8ݡC�{�1�X֋ȗ���zH�<�����#�Sa;�@\��9�ϰ�KKK:[��Ԭ���4��z�E_�%&���=rA����pY �{	m��2�f���\�8#�W���%ڊW�@��2��"�~�j���Qu 6%O����L�{�%��P<_&S0�8{�5��7�l �Z���P�̞O3ZH�ْG��<�Ѷl�����V�	d%����@�؃���e�n�T+|4��X�)F�{���Sw8��Д��Ϥ��������,��x�Xᙙ����N�������� <�l�
�Ľ8p ?��hY�Oa��:�����ڦ�u�H��I��n�k41!nīl�c,r�9��{�7��g(9FZRΒ"���`���HS�o�Z�eZ;$�;e6G��}���8�4fV)��[�C�W1�BS�v�ХL�G�=~��50�T����;\m/��o�mt�g��y���{\O�N��E�b�N�z�'�7V��סB�7~����RI�1'r��2lp�u�º��$�������z��U�2�~�:;i��ʆ�?G8�{ʌJQ��·���@���Q�s�=����u���Ed#ŀ�yF��� ^:�˂Б�!؈w��g�Bǌ�asҧ����p�,/�R������y�&"ޠ(؊��{���(���3ss'vl���׭�n֏<c�Y@sm�3n���FB�[BқC~ܱV�ѐ�
#�e0��c�L�Nͫ�q�0��E�$Q����݅�3G��t�x�8l�W�^��\�RHI��d�zm�JZo�A�ٌ:;���`0�YE]J��:�g�p<9;T�i!����]m4�4�t��������ӊ0�;�� �	
��,I�G5F�$��G�(�Y�؛� Nv�"~MQ���q����l�4n6jfL��c��{f�83�M�ƙ]&�d'�lX�O�^ggseU�=�1��n��O�9u���v�	7��h��6Cd}
��9R�+���+O��]�b8{�eTh/�//4��4�p�[ē����F��d��j��Мwy&�4�Yy���|��͋5�{��ŋ'��S�2вc<�ui���!�C�;�&�n���n�;WgTk�j�à��oA�b�q���MG3�9$"��k�~M���G�J�j\΢�ԡC3@�NwQE����oTtI����f�y�&�x���g��զ��w�kS���3Aώ��1��m�y���tU<ç6;;K,��K�.�3d�&��e���[�vԹ�5�@�a�%i�C_��=�c��i6Q���$c�3k��a6Ǉ2D�� ��#��+Q/+9��iH�Д�l!'���+Q�'f�]@�9������ �>ܛ����_����6	��(	��x
삣�*6��2,t ��`�"Y�DҎ�I4A�i��i�[�F�rx��?�Z�ܫ�������AX >�m�\��!B���)�3S�q��[b�p�8 D.�B��3��Gա�X���P���kx��x��A˄�by�>)�_:��>a�%�V��v��e'R��Ya�)�{3��3Q�b��B��`(Ɏ����RJ����0��Y��[6G�����Uu�2�;��e�lK�.�Q+M�懹&��|�2쩋#���kN1l:��+�ߨ☿��TеV����&�9)�K`DK%
�S��]3�vM���~_YIi8�N����/�����o��� G
��bJ�B䔦	Sњ��1 A�=z���~mmK�[��[����H���Vɔ��~*��!�<�J!D۟�������2ȇ|Q	C�;v����G�w�}����G���o��0�Ӂ欕�@0sss��%%,��C�h���W.^|���YwQθ����p�Y��f��8L?��u����&�!��~-���r�a]���Y�����E.��QU�2�t�Y�N<��J�eW���A����-�}q�r�����lf�z�=77�wv�ᯆa�֭[Ѥ�K	��0�D���1 �nw�5�|��y:��{�o-�L��3�#$��N�{ϝ�lժ�����n/�g���Я0�
�Vm�L�a d+�:�Ν;x�����r,�Z�cI�{����r�GF]��!{�+l����,��¡C��D^��_��EN�GQ�[y�������@���������Zb��'�q���㓓��~w����h�@63��ؖi�v��܂Wnَ���I�A��#h^�v[c�f;���a��J�GIa�����B�U%G(P��vpG����|خo�3���ؖ1�Q���{v:�p�ol��Ȁ�"�B�v�nw�m��]W�3ȷ�8��Ik�F�Y��<�)�dy1�`x8�}�|��D$�S��e3طo�$F�cel�6�����,"�g�+��q��2�R�J$��r @M�\$S��	`"�%#�uffn7�1޼��[���"Ч������_�vt��$�®����<��8/\X,ԉ'�a�~Ig��_�Ɖ�I��7�|��/��tL*/����7ty�*9�h����e+���.�*�]R:ִ��3 �⪒+�ֈ0'���?l�(A�b��OJ���}Q�Bz9D�,..�g�A�������ƙ��\�~E#��q���������{lr|J�-�����w�����;��j�%��,oH�>�g��Qh���K�g�QR�*�(�x)\��71VG����n�Zmd)$�N�ԓT�o� ���2fag��ޔ.�(#��E��ss03�ϟ��Ċ�*�z�m`Į%H�"����.s��\��L	��q�G��R&�k:�܌r%��Y�ͶЯ��
����L-�p�_��0���Q���^�҉~�<���?��a�,oB�<,'BJ�ZB ;���=�ف7$��#�3�m��Dr��-�B�T��7�Y��W&��ǔ���`�
�b�J��sQ�/��h�!�.�T,���0����ʧ��4
C;��<)����l���c9���Y����_	��ml�'8�m�P�5�&M��nF������������u�:l�T�D������O�Ӿ?$���X�g����K�)�
ރM��;��7�`Z�z��3�t/?���ա�Y^O-w�2r��;�o�*��W^��Iꨔ���{�|;L:�Or8�ʀ���0==��p(�ȣJ,��<,�ƅb��ٹ�����[��(�-����[�z���a*��e���6[�F��Bڻ5�.ޑ!G�5eB�;��E�V��,��
��P~�#ݪ��� ���ꈚ�Ӎ�Zܨz�"�vVoWS7�bZN�r�^�\��<?pZI�Cp]-����
���vw�Cj�5?J��+�����۝���;�w���j�%!��~��j���I��A��c�Ǿ[8B���^�y�:�K����'\�4��mq���p`Z�9l�L�BI���b6i��HfN�E�S�YBdz��n�4�(#�u���S�c�䓪HT�<U�kYyX����[�[3=1	g2�QC��L�߼:�!fM���I���s����a�IL��b`@΄�(��ὐ�n'ZZ\������_�&����R��v=طgO�V=#<~i~�/�GhX�sL���<��gfV�<`� W]&�'��x�#8�@@켰�_ޒ�?�K��p�4BdR���gC�q�}+Gmyyu�����]f��Z�==x~wc�FQ��B�Z.1����	�8��i3�/�8]ԛf�R�+��Zz勣C�r�jy:yZ`��J
P)3ޖ[��7���[���+�j���Y���!e�d�$Ɇ�qX8$�����M��t4���A�j�L��A�%�K��09�ǉx����p#X��\��0+�5�m�0�:ZT{�I���ML93wΆZ���-`�9QE�h�2�`���XP�,;�or,1Ke�XB�����Ӈ�;�]�������M��p��K�C�6�lDd���+t��wg�J��`1�N�d�[R�5)I!򄿅߈�5��	��[�)O�����-�?����F&�gB\D>�zS��d=�ߓ����\O�Åi����
��P��%�9F��Nz�֤M�s��駟>{���~�3&)h�hi������^�+L������A�j��BP���*����+�fb��4�Dffq�\�%#��v�wF͇�i@��dP��]¦Z���'`O�$H(n{.��A���t��B�<��p�Ox�y�G*&kMdrw�i���jk��؆�5?\.�*NX=Q]@�G���LX�=�e����@�-�1x�qu���
4}��e0��#���w�dbeܼ���	ڻw?>������&{G��	B�p���e������㧰ߩ����?~����~��� ,����[T&��J�ɾ�,D���q�R�ӣ�"f���<�c�#�������0�����;P�4�w��'���D�Yf.H�D��A]�]LH&	�X���`��$WVV��C���M�O��?�
T�nA�Le 0�<1�KE�!,�j�`^	��R����_���4N|7�r+�C`�L��q����V�����j�z3b�U7����繕F�m%��� �T\҂���"�$r�,j4a2.fDXO�!��
�Z<B>��E�H��w�P�Z��p�&��66R�V���d ��U�H�j�eD[�`x9;��׏�Z5p
cwD���7]I�x��`��C��V�{�L��zS\	�ƋC�^�֓� �2��N��EY��SR��{��g�J���%p��܊di]�=�18e>��̔-]�Cb\ұc�{�q���$Ƈ9���PE����~_��6�����������C�omll��j;Iz]y���/�Gh�Lf��kC؉�"W��8k>����w|���Mz�I ��_XZ�6t�\�E�F��_���gf��SG���� S��6�(휃D���H�ޢ�`O"�F��P�P�l�g5��;�̉R$X�%..	a��5W�w&-:�hz�^��@Lf@�'����.�tB\�Q�'l����4<#�U,h`ep��H��s�-nF�^& �%�DZ9��K�	�C+���пW��~!g8j�5� uz���Vj#�r6���i�^gC�3V�?{����l��_Ŝ�/�5%R����t�Yb��_D�Kٴ�&�	��hY}M��X��D)� };����C������$J��**]��P�8�7�2��i�H!��J��xgK
V�z�񽴐uH��·�th/͕�8�-�K�ó_i�mF52�BF�=��U��2�\�)#|��Eb�mhT4�7�9�U�B�����\�x����˗q;t��
��SH��R��P�V�\�����LC���,�`��a%>ƿ0^{��̏�}/��+c,�C�7r����Qs�8zX�2R�]�Y�+X�Aa�H˦�1�J��i���	���u�Y1Y��ܡ�a�s�{�q]nC"ٴ�7���uf.�����	)|�u���Y��˭}� �:G}�GB
^բ�Ì���7��NB���m�j%ģD !/�L�������Dl|O��A����B8��'X��aW����f�ɌzPw�R7K���X�:S���M�2n?B��.�b�5G���ݾ}�%�V��T�eʄ2sC�p,�+�6Ct/��y�Q��=ZZ6W@�B��O9Q�n�7��>����X�>�0|���ļA�Q�I;�2�E ��Y�U젚J^.|�`������U������Ν�u�B�a�� {����x��x{B�ORl��/-���%Yh�T�4a��:9�;�4kGx���[����37�[�h������f�jO`����s�ޜ�|����$���8�:��f����؞ԟ�� �Y*�8�����&�s���P���ʲ(�v�}����-�K[��}s3ӓK�`�7��2wv9�fE�|���u���r�D�EV����at ���I��V�b���	J�a\����4j���v6{ay�򚝛{��s���ϳ�\�L��������zMTO����>����_���Vg{0>�ℍ����no���~�!�6����&)���"G\��a7C��6�y"S������+��8�>	i>2LS�n�j<8���O�<�gϜT$313�K�[��穤�R�����Z�Zd����[�54*��2��=�g�]��]E��]�(���<���Q����m-���7�Ƨ���0��鵳�D��=:��C#:Ͱ:,����*Dt���^�}%]5�0	��,��2�4o_	�n��/+׬���ږi��y"����_ă�=����������_%�S>�[4?,�0�R^�+��{TO���!]�r<���)��,��ؠ_�r�1b�\�g:k��Εъ"�FKX^��!ǰPZ������a>Le�e(�]�Ae��:�P��I�t��jX�aŰl}��8yB2�hdS����ē�V.š4�C��9�m�1�#�#Ǖ0�@-�l��ބ�,l75�0S�l�g��bƝ�<#8U��S��9r��Mȭ2y��ß�|�6��e�Q�x�D�����Ry��.��L�~�z��Ya�wdF���x�]^���XS|bCC�U�����j8sbY�hT�n"�A�
��jnwv��T
k�zS.K���)9�m l�L3ĖM�f�JGSr������T.�G�LU��Y� �qdJ��DI��X�����n���ϲ�jYO�ٳ���[�n�5W�z��Ϊ�j�/��>z�Ȯ��G�����ReD���qݙ�=��5f1����5�р!e�%���R�,6�<����8�f�YX��q����O���C\�x�'R��r����9�5�Ն���m��`ϟ���=�^Ax��/_�&eF��C���i\��$��l��!�q�9��x���)�+HêW��t]���ݞl�z�
��%���2�W��]c6A���N��R��k��y�거�@��
:v^
,`�4��ړ� �OM�;p`?��������7;;�pdsa�re����:|q�c�8������a��|W9s�U��Yș����]8���n����'O9|�|��F���C���厼�v+p�����^kcm�U�z�{gj8d�%q�Xa.͞qX�(�,�7�A�R�R�I�B\c���ہ[>��c�m�*c�C����{�r5���⟢���� @��Џ�Di��,3���e �pt	.[z Z@���/P�=�Lb[,iPu�y�#I)�)�uIҬ7�?�����\@�V�n7
����L̨�m�[3~ՔҲNgkk{c���?r�Tw�}�����Kׯ�z��k�/�>H���qP{e=����J�����C@4�@"f�y<]��6�ճ�D�I=裾��L����v� $�V�����+W�t#�S�z��l�����ʹ��jE;���~�"�t:��,��x�#��g�'�y6ӳD��%H�PD;�ɯ�A{����,��q��S��lc�}"ߴ�Mǵ�0�Gxw�B�v�ЎQ[��/`��a�p�w��A���lH��}�w��{b��ɓ�>�q4�F���+�`��謳e�h7?VQX� a�877���ϔ�S>���Y��'\'��N'���L�h]1�y���BYV�*�X������~KKK��+�R�����Q�Zh���t}x���ժ����i�3]y�vtI&A\���7�:ŃTL�Ζ�a�;l���ʄ�p��1�g�������[��H��޽�%?�Is�Ȋ��{�7J�"s�!m�L��mc?��4RZN���ڷ?�����a���%В9B��5�^K��(W�L쇕�t�A���Ñbj�ø~��6\ãG�^�zk�/rM9#�?q�"��H��s̖��Q񔫎:�X���l�
@b"�N*�DW!v�UG N�zS��]�3�o�3V�nv���e)��* :�gG����V��,ɯ��A$������ZJ¦��ߴ6˂�"�'a�3*�2�,{�zA<�$�d�/�U���6]a	Q�J�0��'pߪ�3ן�� �w��b�J��(F)�������Ȯ�����Cc��΃��$=�T�%{IlX�&�D666��cX���N�ӕ��r��^��"	�&ND�h�PL������~�H�+�J�֑qf>��_Y^^���d>ZGf�O9/�G�*+#ʹ�H��"Ȗ
�I<���?�����؆�z׮]S�$R�1�V$3C�r0�suF¬�@�Kw�0�l��┦�ܛ��j	�������f>iN5�+����`w�P�>p�.[��a�Z�-ޜ:u�ܹs��{�]�p:jHQ��L to<�<bI_�����x�t�d�2_�m}ۮ��D��rò�&b�~o�Vi��i�:�NC��xƉ7CS�wm�9/7�&��1nY�
�NV:�5�V�`�܁��D'�t�9B�x�ꞅ�fe����]h�w��;4*Aު[��++w+N=�4z��H$9�d�Q.�7'�:��:9Qk�
۳���z�fݫU����]!�X&K��}����ӎCV����R��A�\Aj�m��8�+Pa��&:T�2�q{ �������f/I�A����x��-����C�U'+�N��C?pp_�]�O+�#qc�� �!a��E�f��l��vt2�M�ciR�{i�ROW�[7�^�v����^���Ow��c8ۯ���~��f��nh�P]"h��^h��8���.ԙ�w�K4dA��{�HI�	o#�'�f�'!�G��	��y�D������wMsBN�0�X{�`�=�ِ)Ϋ[}3/,�96�t����4�A2�����C1t�{���T 
�t�;D���Ze�U���XV�:���9$�;�נʰD7�N?��hc��@�1FM8&l*�
zՂ7Dr�"��ŧݷ�a�rvS��v��&�[���[e�fأͣ$;��<�쳧O��NOO�����'?!/���O��D��3���!�|� ��Ϟ=Kln���믿�:۩�\'��� �:�������d�����e���8܈a�{iL��>���#,�~�,'{"�bW��ds&��Nי�F�<�\>����>cN���B���$���Y�N��Xx����P~�Z���ĥ��*����H��d�Mɡ�rf�r��J�l�^�F[gVz'3+p$5�'�WV�z���n����-��N5��I��T��!G61'��"�B"ZI��y�X^x*x�����:bq�8��3g�H�Hwq���'�|K� JQ�X,��������#�] �ru�T�|�	�2#n�<�����u
����|L�*��̺m����S�P�0F�QȚ��)7�ߊ�Q?�g�������=lG�K�R�ܧQ��v5RO��]<��ӂ⋅V�LV���I���b��-����W��z�l��SV�:e�Ӟ=��W0��b|�v�U~��J��������K�Nª��!�l.9���A��d�bTU3d�Xl"qڼ��U2@`�!$�nb��噐�Y8ǉ+��Zm�W���3QES��.���HwPᠴY823�>)�ҕ'�fNq�d��}����B�A���X�e���1ؘʡ�؃�׷�p��5����_�B�t���&r2�������g񙧟~����q^~�e�.8�r����Ț�L03ժ?���.3�a`�N��YP�AM4s�V��P�Ez��^��t���7�`�^���F����<3�p���P��Aݮ��/:bcm��3h�A %�~�J:�=ӱ�;VUx��L�P����-�̍h�O��^�����˼J��%����v3�ٱC�feV+˶�|g��{��"�r��J��#��b8R���@HJX$�+#�5m��m�P>g��c��Fq�:C^�*u~R�k�v�jzOc�a�����g++۷�.��.���I<8�wv�ȡCx�p'��k&��n@� u�u�2�p�8�h[p7����`a�'����a��!�J���8	-��W'���Nrv�?g~�6��=
F�,	~s�)�����؃{�����e�I�b���z�9	}���y�p
�{a�'��2��rۥf�)��>t�����^��Lǔ6LkL�+�D+?��ƍGH�ˎO�Hi%7YVK8֍����A�qRZ�XD����6�s�6c������[�ѕ���2m8aގ�����EV��U�	^�x�䚻v�n��(�)�;4��h��D����zp|�I{a�������|�����a�H���3�W����8�ɓ'���E�82��J��v8��M�g���.�7~��7� h�6D%Im��3��8�y`��0g){����:.g|饗X��a�
�{�SɋzBFqa��"RrpP����7p�t15C���Tt��d!g������t���^o4&���M���Z&� ��)��\{
S�q�*�Ų����r� x
{�h�f�\�}'�\_��^.���	�ٻ�+��ز�,��K��W�L60���b�!���`�S���<q���Ç�u�[C���@�Ӎf�����t�����m��	e�Pw����FC��C��R^.RN�6���Rf�8\d�T�4�uy��S���V�Va��$�_:zI� G�d�<����"f��d�o�(��V^�5����2w�f[��D��8k����G�檒$�V���ZL�h>�{A���!L�|�? û�4��r��<�ֵ>0H(k�- �qCE<{�i|�-jxP$0�2���>�9��I�{&�Ҭ���oWB�B���0&�������c1[M�����ȸ/(4|�СC��){j����@T�������/%�W�����iIG����r�k�*sX��Q����}�#h�&''�3M�˸�S�N���H�I�Z���A��p*��ހRY�n?s�x��]��+}@w�Y�aw�ѣGanp�?��O/]������ir�pӠWH$l��O�<�u�7v6�l�O��0��l��+kи�m߉�d @L�
j��h�y}b̮7�a/,mm�Ca_��dI>(�ȱ|/��5Ʊϭ\�kIԍ�w������l�A�xy��k?�_����"��W�v6V�"?~h�S�?={�ɻ��jo��d;���+r7Z�	-�Xv?@<���z8��[a���j�}�ȉJ����f��|�4��t�v��<�F�M�����ɘ�����Y#\�eR�	��hǣ6ʄh�Ѵ����=h���5es�ӟ~�WN�8Yo������O~�յV��on�s�>���O�:u
��߉:���a|�%y��]�����T��pG������i�L@^�.�)x"��}�6�C�����ʕ+8&�և�%��	@��fkq��X�t���J��y^A���cI>DPY�r/}�|��a���C�*:��=)zӠ���&3�̓cc��;���Z�SԞi5����d�cE����0���g��ؕf����Ϋ�o��a�'A�0�rgZN)����KW��f�X3�0t�Ӝ��Z_�Uonn«`G�ٱi���HN�$���e�;����ϳ1]g8�׉��6�������@@)���Gr��1MB�-����D��7n���3Ĕ�/^D� �1�m�`&����Q
�1��٨�S?��8y/��[�1jn��%�������ի���\X�'�|rff��r$��0a�r8L�88��8��� {���<V �)�_�W^A$�ۿ�۸�o}�[��ϐ�J5��DQrħ��~�*L~'��>�
�>���'������j���I���u���0�eIg�1��z����8�zy"��x��cS���f�빙e��¦:��l���2)�#*2c(I�/aml
���O��رc�<>�-�}���.Ćl�[� NN�� LQSp�|` T�|��恭D��|�}M���|��@^�>)��5�M��h.
���Y�^y��i���h9�ӆ@�N4"�<,�����m��)9���6�rEH�4���G���ɲ����y��
P�d�#sD	��I����6s�Ҵ��x[#�h�,bA���hF�]�vZݍPȇ3��7���*�
{��n�4��lXUx,�suu���x|���^W���-Yaم' '�(/�Tk��{�'�6b�#lR�2�t��(ae�+ɨ�ʕL����r4v�v���
�e�큍U��WI�H�<z1��7���?��f!?Х��r̩@NY��
�R�t�	K��/��_'E>���E\m*�4��%��t�{�_�����Q+�Bfr��9r䳟�,��w���[��p�(��}Mw���@#�(R!
*�)7K��ׯ]��0u&��ث��t�I�S�m?-�������Ǟ>����w�ݹx����X����l-�՛�J}��Z��?�������������jerzfbr
��25Z����SzV���ƍ[w���0�JQw�������~�������ݙ��v�51>w��(�#_�Ri���fƢL��2��Dn%˦f'NN{�0�
#��.�qBΜ���:MLá���� v���y5z��Z�6c�S��I��Z���LE׸x��ڹԷ^�>v����=����^7�������_} Ӝ\�8v� ��nw���+`�
\����\q[�UD��e~emmzzQ�0��u��`v��J&��`���-!oߺ5�'��k�w����g��ׯ_�O���!���z��	�C����Z���D�z���S�	?cճ���!���\ő���9�?�Wq�3<�p����i�a_�@��"Yzv<c�}�
Ѯ�k��o���F%�Pb�+�v����X+h'Y��J�C-��ҩA����?�4?�鉅Ss˨F�s�Wгd�Rf��������|h�V��$�V<7c%�����t"L�b�'��lN3��]���;w�TE�TBp(�5�qL�|���'�+Tu���P�k��pm���C��G�5�	��[__GhA��hAqp���r����+��>�|�Tv��a�/Љ��qI?��Oq���z
������+�!����F����D�S��Ν�����9�]���OhF\*�1.�m	�zƣ�A�o  8[���h/���-��8������� p��k�"1J<-��h�s�E�Eˌ5����9�Dw!9ו�u��������>���/��?�����6�8*�8	m3h�qv% 9�D1za�U��,�ʅq�x�uok����1 ���0��a����nTeu�8�)4�ܭv��k�I���mȝ�zCv�&�BE1��'ld	�ϑ��_<&v�A KZQ�b�Xq�3�̐���b�,^�HMo+�M�k&�z��J͏pGཐ������k7�GI�`
f�V�pj�����U�u���l��%���TZ�&#a�H$q(������!�$\*En��&k>� ���%�A���u A��V8&��d@�Ȑ	o�ۡ^�n��;��&�l��-���Z����L�L֨�T���,��4� H�x2$�0�0XC�R�3/�'��i$�2 n:�s�eb9mg�SfY�cef��L�]p���_�B���?�z�_��/���������յ?����Y����ɚ9v Y�r
�<��i����n'��	���C��z׮\Y]^���p0�X�''!
������ع���w�0�|)���>,�������K0����>�z�T1��犖����h�_�X*]�M��ߟ:u
���ŋP� ��4$SH4�,'�����f��3��DGXXX�m�UY�&&�h��	'_��={���/]z�ҥKԜZQ|�OR�~(�>��Q1V�{_z�g�9�k��O_5���PzU�d�o�;JEG�ȝ-l:��	�ߥ��z�׽��XYv����fiwuu^��n������o�����?{���jq5\��j�9�t�>�LQm֚����]����Z��v��[?���omlo�5�}���^�5Q��NV\��w�����Ûa�����u���Wݢg����?}�_�7���F�7��^���[vo����Ǟ~"m�i���H�\3IF�R����y�;v?��w����N��f�Kwn"��"R�.����#���U����<�Ii�#�7p+X��������')����2�r'6LQ�p��.Z�:"�t���بՙ���VD){n�g	@/����o-,މ����ퟶ��ࡣ�nx�ւЦ"���+�/�<�|e=Ы��:�w���,� 7�*P�ބ;6$��Aߎ��W������p����=�(<������*��^C��s�=�"D�WNW���i�܎/��]XPҗE=�G	6Q��!�ȭO^	��A�L29j&��p� vR���.�[�a�%'㝎:gҢ<�MSS��ZT�{�W��a����q�s�FMK�Q����Wƺ��X�aXE{L6X�yh �套/mcc�'2Ma�
�W�Z&<�+@.f��L5Ɵ&��R33�Ӕ-�.Z}�	��&K^lg���i����"m|b�
AG�i�wAT^y��5)>kR�2m}b�`3��iW�h'��_'�idH�@u/��&�*`8��N��zv"�ʔAR�0I_|wę�p�<��I��p�|v�k"yxdkgI�_�h�Z�)u�xS4���a&��A).��SzT�����a0Өl�bN\)�2�31�CF�"�pG�0Bx��SO����a�})��qĥW�����H]!:Q!L�i���f�홞�����:�`��M���~̤tQ8E^k�{��3KMWU�p�7�����Ic�d�-Q�ٳg��x��#��G��7|��A���OЁc揌��,W��'��㌸B8�̀p�Y#r��V��Z. ��q�Ґ�v�}3�Nn�jeZ��o��
����4z��{����:�eTJ:"�����D#��yX{Ҧ�9�yX�w4��JE���g�ݘa�"��b�Xb�N�ś�(��F��;���嚁��'I��ֲ����)���J���1��-�ѥ��T5q�+W� �k7�!�_�XY}�'?��W����|�N�>-��V�t�����Tk����(�]��/_�|��<�եKW�~�]]w����w~�w���������cJ�8Y�=0��}A��<#^�U*���ϲ�,_�"�U�y@6�3 c:���W�WP�:�b���<����n�F�a��{#a&"�W^y����2�Oy �$���r�1�Vj�Gt�	8X��/���p����˷�z�<.�eSJ@ �����P

��]3����[U8��a�Y�<���>�ę��6��)�p���#�=w����־��� L��c�Mlx�i�Б�pM���w�^��ڜ5�i�J�~8����NH��Ud��W����iD������Ӟ��յM�S�U�zC��1E"�������N��ٺ�����-��jV�0�LS�kee�2�a� tא��É4қR�x�n�ڵFc�*��I���"���뛣�X� �"Y`�a�1� �s3|uu ګE;2OfM�1	>��_�⯾�� H���04���0���۽nn�WP�LNMq;�2�W4����kbma�����(KX4����Y�B��y�jl"*6Q��pc�DǏp t?�V���k�dA	��4�+�vϨu���K��'!�G~)xI9����`��@'��ԃ��g��j�e�s7���fC�>��U��h���XEx���`,�(B���'�0㯬6��&r{�O����@�����J1�Y<P5h0��o�X�Pb�2��R�1b*N�AK�#��d顷A���f$��:��=��?�[0<��fSk
V�;9����fT31��,$:NǪ0	��e^0���J�ߔ��pDe���e#V�xsM��b!�%�˯]���;�@9r>,���*���0��� R���5�(�:E�$9��+ϒ��`Ĥ)�^�T�.�|�����^SN�Ê�p����Lc�@��6�M�-�#�n4i��u�=�w�]��Hֶ����j��kMnow��'�ϫ�ăO}������f�;���ٽ�%b�����v�8lÒ7�㻺���ܼy��y����F��w�5��Iw�ر��{�uW��g^x�L�C��=���-F�6|G�}���\�8>9|��4�(ŝ��,Pf"Q��2^n�W^E�O
�J�s\g�ը����F*74��O���1�~E��@
Ω�e���ް�k;���O�⤼�e�e�i�H���URY�T�Q�Y��aI�wǖ3^*#2�'���^R�m���5m�LN��5��6�����*�`₳C�<��Ä@�}������-�}ǔ�_����������������&&�{ͭ~������Ƹx��$)��y�������ܔ������7�j�olleyv�ԩ���o���B�4rxtW�S�7��|�
u�
S��P$-��WA�Y �|���^�n�O���d�K�&�`y�9OD�-׻xa�n�µa�#8$����:+�J��Cc�
ѡ�:;E��A�ˣ9��Jg�����rYg�>��cg����^cF�8Oe�+�@	�lC�bëܑ,����q.��Dy�7Ps1L �1�,�_k��Q��f7m5'�aRd�e@��Ka�yf�2�2E$$�$�__����^y�/��?�ez¤�������͎5�B�,Lp����{o��Ϳ���p�ƍ��������f��ۊ��6�V�cu\Q���Ezsǳ���P>��~*�5ZY�t#��˵2��0����<��#���c$���+�z����ɟ�	l����'Ƨ��F$���O�<	�_�ט=`d��BCVLK��Is���~%h��r�c�����9� ���]~튋JиQ����k2���e:�%ʌS[F�a�v\�6)�K�IniV&+>"�ѣ ���QU���	酨r?1)P%�0vhVbl���Z�Q�E�Iy���,�Pf��ᨷ������[I[�����B>ez`4���ׇ'_�pNt�gT 5'ʤ,��hV��2�yV�X!%���,Vi|���g��9�m�d�j�2%m\F��A��J��>:C,B���K3�D *ø��7�t^k����*��d�L!�q�z�&9�'�)�-��b�ÁnLLҜӥc��7�+��Co�&"�.��
ɞGϘ�Jy&�ca�?���W�c�Y�S��O�����\(��7�'k;��K.\x��g~������
,z��3hO��g��X°,TȾ{`ﾣG�on�dIب�3cRd�or�vpn,���붋�?{����>�+w�o����2;ujvv�,�k��������A�����0��{f�k����xȲ[�1n�믿�KE,�^5�<�!l.,#=6���5D�F�]�X0�ǳ�A�A����(��c�īW���a]�:&���$��e8�uA�[�M~�̑U�|ʠ&kD����2>9�c�\Z�ԫ9w�w#|��|X�aP����D�,�TG�i�&,ԟf����"nİ�%}F�l���`��#���TN��\�Q�"�ðG�$��Y����qL��h���a*B�f��3b�:7i�M�r�������c�fP��򲰴D�W��À�ϙ9����0��A��)�!���]�z������ �xj�$����������(S�[��P�\�R��L�Ѹ%p�C��u�����:�G�x�ô�ٳgq��h.in�MP�2}E��H�\������2��1,�s��ئ1��?�,���(=+c |�����g�"
�q���
�*H�b|~kD�6��d���Dy� 	��5�Upk��e�S��;�ci�D�t�w�{Ǧ�[[�~/������GVP��HM�Hm�,/I�A�9����EZq��_��'����_�t�K�g�܁ߨכVа�Xgl@i�zU�W._���O,t�n\��:�F06�۾�k�����a�Wg������1��"�la*�-A�s��trgIɊ{�UnM��Qr"l�7�;�0e�n5��W����6�����GLL�?��>��O��ޢ/C6�@t����L���u�b���>}�	M�GQO�+��h4�0��N?&e���Ux����n]�r��5��#��M�'ˆ_qG���(�A��B�I�*UG/Vu�)���#�q��١��?>�"����aF�;�6l'���X��l�h�ƕrΌ��&�H�`��$�>v�2�)����/l��Z�
ж%���]YYa+.��y;���ƃ�B��!���R�H��ᯰ�Gr�"��HL�:�o�V�U��_�W�.,�[xFXp��.\�g��Np��b\3�"��ND�qbC8V�X��a��=z��Ʒ8��c����_�:p;��'NU�ƍpI��#f��H:�H�
�MI���"��t�,D&��"�Qd^������d�9��WJ.s��"���Ҩ�2�.�X!��dRj4��;�"Kk��۹�8�3��NK�@�p��N�=ْ� la���9r�/��W�Je߾�#zɭ����]��qm�B�ׇ[����X7`���]y�ҥ�>|��54�3x�x��ʝR�
�^HW�u#X7.��⊿��i���요z��z��V0� ��\@MWC [�L�p�(��=��$M.� x���a��~d�Z���k��@a��Z�U%�y^6��^ѿZ��S"
�f�b�����	L"��>d�ȇ�7ʨI'�5�b"eAtK/��(ZO	o$@���J&��B������e�S�`ֹ���ɉ�$��[�Pm��,,,3'B�G����`)�x�Nu��!Z�n��`X%0iAڎ���*2�a��!�!�������beh���NcW��=�7'O��慶�ffOSK��{���19AUk�jθ2���#^˿C�Q�tD�{�HȺ� n�(�p��ܹs��������[$C>V���0�#O&���b!9g�<z��7o�_�g5._����a#�Q����Ҹ�@M'n2i��2�h�'}�d��Xu+���ss��y�ٽs�p���1_��@���q^�P��-(f7��p'�������d�^x�	+UN�8
�왱�Ĳ�"��ev�݁u�¢�"\�YT�J%���y[�n�����a,kH��U1+�:�a��v��)AgB�>}��	��#33���|---�b�~h �yA��D�flEB�1�a\�+0��D?vM{����܏���?��V�Yg&?�3��JM#�I�Q��iF��7�|���h�S��/�.�uX5�����:�6A*�#ٜ�z2��I�a�����)���'��/N����(�Cj�`8�ݽ{W�YG$�d�L�+���R�[(�?�W�~\��d��?���p%�����l`}饗`$`��|~����������)w%�!���Xgr:kjP���j���W.8}_��/��O�K&�����4!vݺu�#e٠�tU��z
?YMRj/���+�:[qpXh|�^���X�;�08>���DأLQdԧ��=WrF�dA����B�%q�|O)eɑ���q�r�P�2�80������S�-![�;�D�L�Y��{�^���ٙ4�<~����~o'NB�s�
���T;ʊz}���Zi4ܜ9s�{�~�'��:w���G�H��~wǴ�I@%��0~��Z��}iJ"�P���/{o,�y�	~{�w��[�^%�$�%k1�j,l�n���00�LL�����1&&`:�����nh�f��X��-ɒJU��T�r��Rwϼ���s�'�O�$ٖ-�8�V��f~�-�r�y��&��R&=���h{Sh�E2��ֺ8Õ+W�/���qu�Y�{1���9-�m5�ww�O֩'ɗ�}Fi�(=����tؗ`�����$�M�����X�^d�̹��x0��벡��Q�f�PRz&x�ކQV�-B�p�� U
�67u�Wz4Ţ�&e��9x8@h�hd�0x2b��\��эH�(�!��.-�xZ�t���M<Ώ5�*MfQ~�g[Dh�績�	l������V��F�k׮����(Oh�k	�K�#��������J-��8NY:>=���ů���ö%t�׀$Y��T񀰛(�JoO��m��z$s+��u�-��o	ق�v���>�n�7��yft���<X���5HWx�Ki��ՓNQN6�ң�$ux�U�.��za������o\�����u\_%��;�cV�lA�A��#K3���T�n�پmz�1�Y��������.�M�H�#�\�R5�M��Oy�6���vӓf�F&-�i�~�&>��re��|���e��4t���i�$EO`�t3iѹ͎�(��Mמ�������N.ܮ�+��/��^ݪ��فASH Ty�kKAg\�qΚm���������T�f���m��c�����R���0�s.6u�8��sӪA4��
���q��du��A*�ۿ��Bo�ֲz;�ױ[�2���	ya����K;I�E��5[|�z��N�HJU* &_�Zm�AVHf;*�ܹs��XY%S_���U�(Ѣ?�:����ur�����ٌ��0�Y�	�9ˠS7aO9u�R�.[&�q��H 
�l`�bS���/m���R�,�a�[�������\�:)i]�Tl���5|:�k�� ��� * ���@Ò �6l}X��>��l��5�7U >g0-�_iri��ƭ3"�2`zg��_�;55�\2C������˗qϔ�T��K`_�t�.C�[�{N�rXH���x��������g�"#Kde8{�,�4:��k��"-,C4Lmg�<��ڤI�I�Y�O���XN�Mk��-Z��N�d�a>���5�۽����%��%S�,�,�1�A�;+|���"�8q�ޑ����l��5|�����������R�lգF-ެTgG$��P��ٽ�o?�w_}�����D�(*o�mm��Ɠm��#��c��i�0I �DU�n�7n`�154:�'�Ƽ㴰KX�L�M����ك��F㜘#,��O���Ho�M��I8D#L�r&�X��2M�z4���Jp��+�z٪��b�Z���Ku;f�<�y��L7A�̠�{�2��:X�E��;�4q:���s�d&3�������h%K	�FŎ&oԭ��Ϟ�h�VJ����ͺ���Ôp7�5�ꓫ���;��Jɶ����?�C���O�y��UR��C�Pu�y���s/c�I.}N��Џ8��\S5B�:����@�~���򗿬(��S3??�я~�������?��@M�s7JFr��@ɧKb�[���V�\�d�]�(���}8�LQ�s]�x����Ld��Uy	�M����Cw<,*f3����˶,�d;�mA3�}�!���
r���gΜYYސ2z1��}��z�_�ޚ�Y:ܕ�'��}�B`�n/)�睶�|
�v��":��mA�onV��ծ ��U��1-�b�������a�Q#�hnsaimy�	�U5c!l���ñ���R�mZf�kQ��bf��=C�;�5��v����ܼ|}����}p��e�;J(��faO�'�-��V��]������P<����d��D�3zo-?{KΧ�;�>�\!l?�����v�U�o��3	��7����$y�
CT]k$w�Ե�n�,�'&�m�M7>x�ח.¡��xeX\CF�Rii𴲸�O yooU�6������|t�B)�c�4t�3��A	�����iN��:�C��![(?t�SF�p*�k4|y?TB�Z��3������'6?��o�J��x:M�+��'��u�o��]ќ�%hg� h�0�������e0xd�J�IB��B�Q �D�f�=��눗�	�R�������ө��D�ͳs+Ld���СCxF|���i����h�R,c�((]������&.��ѕI�ȴ���UG���M���D�|�pi<�X��yǵh-i�U���Dz�
��H� ,Q��?@�z7kk\�\��ǥ�%Cm��Ǐ5�c9�V=㹦��%���H����0(H~]��-�o-̿�����G}�о�~����XZ^�w��l�m犥���my���,�/�I1V��pѮ]�����7k�z6��[-�d��f�j��L*͜7�P�\���
prr�q6����4�V�a�K���W��*����^��b���Ȭ����$��ߥ��|���/M�#.���'���&`�nU�5��v����u�_[e�p�1��7@���][['�ͦҚf�AH�$i��L�?�a�h.�VZ���D~�#HS��=\{؀�Y�"��E��p��)?�N�4�ur��:�2D��l�.�y_Đ³�_�ˤK�%��lx�W*�H���������>661QR��c�ç�~"�LhL\�T.�U1)k+��pZ��~�������/��O<��F�s�w7 	�v"[��L����$G���.�e3�Ax��Kyj�ͶL�$k"U	�k	[����\Oq��S���?'οc���b�H}Q���ن:��;[�m�S|����}������꫊JQ�;����:z��7S�̙	�m����;������5�SH��M������gl`��G`��W%������P����.=V�t�F��k�(n�3+ ,S��,56W�!�HqL`��w��gdS�O��eY�|)7<>���m35b��;w_�x��7O�n��vynxxԖ�
vĝv�;V�qX�l�	̨c��//V6�S33���o+�Sݠ-i'�h��&H�J%�fF*nd��&��4�8��sV�	v_>�5��^�|�����!�뙢0��������������$���hcuՏR�L�IôM��� ����1�x���K�������V�粥�V�5�������͵r��v�!V&�[�,߸q#
��3�v�d#�_mO0�AEK���xtX2�M[������k$�Y��6��X�G�at!�a4�3�ˌ�w̹b�v6�����2�ʕ����'rl�CХSnx����>;��uM-#<\0���U�O��gJlK�*���$ڷo������V�c5s����pH9����]�=F�X��ұ	L��$�*U8N2==�{�n�
,�';3g�,��[|�ߎ���� 1'�a���<y� �Ԫ���^���<��:#ı�?!�dQ1]�LelH��2hC�������Ϟ=���yG��,��%��z��	$�`�x��QWx��Ћ�I�6�|F8�V�T͖L�/��@e&�a`�e�N���J۫啺_��6޼z>����9z��7.�?���*���Y�>�Y��G�v�a�옸��LÊ���(��;vb*_z����G~³�G�lvmsKuَ�i�)/E�N4�;aX�ĉ��ҥKD L�b!�XW�^��ڳg&EW 3@̿r�a���c�=���W���4��&�^i|CzF�݇Wsd�

J�;!3H��Kwڔ9X�[[�n��|���f�sS-��a��߅��b)��t6C�J*1cU�K�����!c��Mt�$�gfK2�M��P���89�3K�p<�B���6bf��,%Wv�R��.)�(�e������[���b& \ުtÕa��(w���B������S|�� �n�%��M���"B�j��n�^��dĀrR�Bq��������'�|M%�"�\��J��������a�a<�Ǟ:��Cs7o�2�Q����X[X�u����o~����UF��c�$S��W��������7�/��i|�92>1�c3�Qm�����?��?��?�c]�IH�$jc�uY\�Xx���L�M��ܶ�Iw�Ķ�t�D�}�RrI�z����O����Y��ꍐTdɓ��mS���o[O��%�F��T�Ka��9v����ƫ�^_^�`]���CEr�FX���R�"\q�9A%|Ea�v-߈���I	Y��vi�eg �-�hpe�kHw�#�8x�#S�o���)��o��z�̙���fwI����Í`K��n1�N�իQe���b�$j-�K�afS�v'0l�P��<LҎAwvr,��[v&�OM�����t��v��/[�KG�/��-�����(�K�B�(�`�s#��w��v�yυ�����0lF�%�l��2UFt����9�5�OI�y�4�w��п8v�^蔫7�^�r���(b���B:�n��A'P����ESW���QU�U�O���L������g(�D�V�n�$�^\B9��["dm&�5��������Zb�Eۤ�.>т{[s��5J�� ԗd@��QRL8���;u�&C�.�3��&�x�̈
��IS��y��J�_���"D�s�4�S�Ҍ��R�d�d1&���g$=�clr
�rǎ�@����:L*c���T���t ���u �_�S���c�T��6E:2�-�3�{�'?w��wrrV`#f��a I:Dj/�j,��͓� �� P���uV�keۂr�� �a����ל�j���d<�9ښ:B���I��r���N/;�c}E��i�B��TFE�B�n]�����<2<FC
٫rR9���]��Sma�R�J����oK�K���x��~��:s��_y#
�����S߻�����_}��g�My�#G� �g�Y���$V����vS�*S��sǎёq���V�Ҍ k##��ՠ�gs����z�r;�$���:�7����%a:�p�/�x��1���d�1$P���/��2�>m���Y����'�@2e`[I��$�9�:"�:����*V>��S{������JH�aу�!��g�ST������Q����x�IG�C����7��s�������-`qr�����q�v1R.����a^JC��dK4W��l�%k%��"��I[�I�N�����/G��o�F'��F�kLLL���!:�	�繹9	1��;��׮_O�2�l��+�.��&��T�-wݍ�&>�:�dF%�p�/!Y�IdS&L�"i3ɓ���HjJ�ID���]��i�-�A2��c5��2�������Z�S>�HQ���=�w�}{����+҃UR�hP�,|��x&��-�Sq����[��B�v����@Ry�*�B6�:i�n֚�Lj|r�Б���b��nz�.�y!9PTv���a�9v��p�0Ei/��g���S��V_i(��Fl��Q�f��>��"qdd��:jX���:�H(��|�������\;��,����z��	�س��;)+��ϴ3�B���l�,�y�=۰����i�8�P����#S�+��j)D�=z��>��ѣ�3��핵z�q�z����Ѫ/�s���ѪS"F��,�*���n��/�*K��d_�x�9$��>��Pz/@k��Z�6\Ƴ�8_YY�9kf|prz�ƭ��\u3.D���zipHO!Q.��dlM�����Zюgm�nF��Qb^>Tl�R`��hۈU.�Ɛ�'�9��C4E���"z�ע;�E�D4�U�4%�t>=!�V�S�h�B�"�	�pζk׮+W�0����,�׋�>-�%�ҨQ�C��B7�ΒOʳNT@cc���.ݝ�>l�5� ��7]~}������㊗.]°�=�⥗^�9�=qT��x�{ՋAZĊ���/s�0A�av:b�]�i��H[	�r&�ހ� X�,�a��kR��#�V�)�4nذ��V�U�4��:���:Vf_.[�a�}<�$����n//]�~g��}]�
�r�T�|�R��a���������F��kW��'�����*����x��{�/?�++kXԩn����V9_H��N�R�'��xr|b��Nǲ�v3�Kg`C��O��
2�:�Îx��:���¼c֘���b��-�8p ���.~rT�0@���֤��h:����|6�Ir�l�B�B$�ph��i��7]$�p�'85������ۆ��ݤ)F��T��;*��kC��UtΕ.w�Mƒ	��j�`��@�	*����m�3���m_�o˓�zv������=���v�n�"�;�e�����b�A-m�=.�����}�6��H�w�O��7�8�M�hW:�Y�`�Hr�B����KyBؠ��$��s���3������\NZ��<)�b��p�Ν;EAt�������C=t���7n�ƻ��L�:p�2g�\���X�dԤ�b܌��p�ד�5Qж��9q��*����ݑ��諾q�ЈWܳ{���,�(2�m�Zm	w����f���([q <!�cib���,��33�n������H��=����>�5��5��z�Ѫ߃�\<�oB�g�����[���ׯ��[��gK����5� 4l/�����f���	�>8=�'j�>����ә�����������t$�as�(����Q��V�ڎB�8�KeU�iZ�\��c�6�=0U��O
y	���ꎬZ�vڏ�6��,�l��=G��{>Ce�Ѭ�`J���fF����Ԍ>0��浴8?>1�u�;�A�	�K\�-B�x݂A�)S*�S�`V�r�$O��>1����]@�WQ�`�C���L@����di�6"D���Z)��Z���_۪�M����Xe�${�׶\�mPL�a�B74	2��i���b�<K��fE5c&8'�aѴe���ę �� ��~�*�����=���̡b�y�i�t�C�.T�`M|H.>���k��ݢ^��F�4� ѕ<IEEJY�B�N"�`t��2�8lll��h�IG�`tT��=��B��k�v���"��|�2 �9v�,~�������b
0;�IӤss�S1�0�!G�n�+�q��<�L���h�04�$�6s�ȭ�g��#��C�6��1F�?�1�/��~���A��d�#`�*��a �(�R�f�^k�J��٠�d&��������;]�/=�@�$w����Z+hbl�2R�.�a?NNN.,,U6��&w�2έ�[�c�s�}�
J=�BM��r�g5AAvZ��[7q]�I#���p��E�(�M���d}��XZ�}������  ��H|cE��}����+�`l��ۇqE,p���^x!I���l6��	�c�_qa'-����u�:��A���ͮq�/�`3�l%��N��NG$w�U�6~#�ʆ�nt������T�U��.]�{����v֔b�<����%u����	V���Q�ђ�l6F�L
?Y����h+�H7�n;�T��BxA%��/�I�;MZ{�Dg�N��w�f������3sX��4$����>77��el{)��,c��/|��W%!#���>���x�y'�ㆇ�U�<���� K���R�I߰f;d�1>�T/C�f�r�$
%C>O��xI��7T.u7�1��A��W�-����K�|�{�5

��Jg��q��>E�#��"��t��j�,,��\���noI�"�Ng�Ŗi�Ό��N:��t���V�#z2^-o�[3�X\^���������͛�.�\TW���Tk*�kņ�[
�t�;RT0n!ipm�'C�t\Y��Y����K�Wn��T�6W+������+��Lڹ�f岨��h��g�fl�!]$F�l�P%�P��nژ�Sa�g��?�#���v�̕���J��~;���V�W��VZv�0��}�Z�^�(m�&�����V��D0ɳ4��{4,Ɲz>3H�ߺ+����/����Z������2�hƘ�R*���l�0ӍF[�y�a�ף0�u��S���M$�iJ�E�iDlC#mt�=*-��	*�oq�T&�NPi�Y����^�JD��i�p�����&�|��ՙkOG$tsmWi{�!��qc�t'�ː�~F�*���"W��m�it���!@ңiv,f��,Z'�Tum�8��}�HT�3+�'n�������333�=/^�t
�)��s��)��^e�0΃�֤�-�f̑���12��s�N�z�y6L1lv�!lHI]�_M���
��s�J�SS��a̍g�?�4�i�����kġפ&Ig�qo.[��b��V�-U}4$h��t�6�	�ȓ���$Ac�Ύ�R�@�Zf��4�Y�:��� �J����W7��/ySR�J_1�^���ɤU9l��MS�m@�NN�GGǌ�ǌ>K���� ,9c�Am1�f����o��~�X�F��tq�cy�8q��+b�Ν;Ǩ#��hP���c%c�Yw��˷���ƅӳ2�`ů饀�qK�z���"5M��q�Y��Τ˵,�ݍ�^��$m1��	qԍi�*� �P���:�N�G]�������_��N����d}J�W��j��V˳D�*��au}�D��dn��Q|����8u'�´�YIGe���H�$��~��m�w�̩�(�ھ/L�v,/�6�>(�+W�=~8F<G����XBl�Ie�:�6k�ߘ*����
��_4�J9�<���(�b����֚��B���������E���q�A8y�P����L����AW �>&�����+++t6qĠ�0��!T�-K�0@��a)����J��p����!��`��c;��n.�eg����V(���
Qv�P�Z>c�;��3��vC��s�X6�
�[$�3RĔa�C0�-��+���y��?w����ά�77�#�"ٰ��<hZf�P�f�q-�S��تl�;�|1W�w`k9+�Y��jw
 �ޠ�ΜɈ���~�5z����Ꙛ��c��;�?�m�Nynzmu������:{(��p���(�~`Fo{AABB��<�8zG D�)٭��6SV��"�>B�礔��=㧻Z
��T�o��0h�3zk>�M��,+Ј��Jb�a���b.?5!��֭Eqr�v��tJ��Z�j�U���Y���+�l2h)� qZ~�a��d���:�m�sx����:�!V�ٳg s��:�GJ����֪jc����S�ΖєJ:���}i�ID�����Vqf�
<�������Dt���`=�N�����N��^��'��o�`��3˸��<�,����<d����^'O���ge<����`��ǟL��W�dݼy�UG��w0���%:ْ���C�/_f�=��h�3L2�\���5�;��~T�lIĬ?�mS��	-"�����
$e��rq�h�>o'ݲ��꬙a�&za*�H�	��-gJ������p{���]�N��!O�;QǏM��������_	�M�p���ق��7�f���s�R�<�M���

upp@Z���[�B.�o�>��t�E��rk�P{��g�	�K��3�ޤ:ց� �w�؁߾��k�hBJC�s;`y��G��Op3�
hW6N6���Ո5Id����;�ak,�^�A�mK�)��Q4�z��h+?ٶR�k��,���D�1������S��"`�;�E�G�B�0�Dr�FL $�28)IJ�.�ر����W�7: ������sņ�yr�uCӎ�-)=y���v�&��kg�ݸ���B� �]M$-�`O�aC��1/����{���=\�M��!�hR3�X_(U#�u>���^�ڵ�!���CPp5b'�A��)F1D8@dA�0�����It�����>�h�����U��,�wi��-�5(�Y��?w��u��AH�����d��Z�-��N,�{��R�t"G���I$��Z�2MCb4fl���ŗ_=��dK��fB�	���u����T�mB�y(v�_7l3�ʹ����6*��ؔX����~[��p!/%-]-��ʤ��*�~��;<��X4��G��U4!�J�ҶJ�|�0F��m1��+��k;z8��k��n���G�Sʽ%���8��PXKa�K�4����{��5:���ھYm�����|6700$�8R-+6? Bw��G���u���n`�kٱsY�%�c�����D�^��;9����v��i9��o0'8&+%a69�c�w�|`�y��U�T��>�m��k�*lK�s;�z�tď��$��G��3����&9Z�4^i��ј�L/�C�E��ih��0=|�05���,$Ƌ�U��$3����-����dD��:ʡK���H�?C:�~�i-��B����?��Ő�Y��>�B4����o��ux4ܕT����fN����-Ѳg��.��J�Z�4p���:tg�5���O����/�J��/�M���� �LvG!38S����K����I_<��X��)�؍�T�l���l��X���ۗ4���ID��	��㜖+J]'�����1�8�h&+�RSS�^W�ʤ���:%���3F˳̶ro3� Y��u��6�V�<7w#�M�{�l!�62}%3�|:�
����Рʗs�R�0<2�q�|����ȱ����Hٮ����Ьe:w���\UF�9}��< X�~��5��3 ��	�;wJ��X��G�t��zboVM���P�]-h���u
��lwڤ�@��775A6Md�=:��ـ�8x�\؂F�;Q�TQh�܁9#i]�ô^]*i$�=b:�W�4y)�ض��4�8Dn�EI�]z!1ŲLf�"��ᄶ�i3j82|x�N��	�cKw��vKv�M�P�.�T�ǰf{�����a�6�¤:�F9��V�N5�0����"oKp5��æa�����K�奥����~i+SHJg����Y�m��'.�^j�xT���l�<lB��V���@k���Å�2���[@�|>8��]�-�D7�.�
�V5Bz0q�����G���4�R��v�i��8D��,�C���3�LlC��i��u3�k�֟�׿�{l��'�ohbwG�o�0�-���\ϖ�9���CA�c#Z)Gj�\ɑ��3��}�C��l�	�J^e MH%p�0@(잖�ڞ���7�S_yqr��}h�0T�%7.�M�!�6D�ӥ�h�.��r�N lzAT*�w�ܱh�UeP(�i�@$��γ�9� �7@�1O	ќ�͙��ɩqȜť�������Ņ��k��Uh������ ���K�D���.�ǘ��K��7V���s0Nfv�y癜�������n@H{Y�t-ǒyƢ$�B?ЬP��=��7���U�p[��^�!;θC�Q��LWXTB�îչ�S*�Y`W	CQ*�3����L?m�j�)=���C�0��ه����C/�>H�Fj��ƯX���&� O3b׮]P9gϞ�q�~k���U���5H#�mn�'�ØT��	��$ˁ���H[9�s�}�$���� ���89lG<)���\�a�1�A�N�Ƈ��5h�l��N��@A��1��$/�@�n9�?�v��L�4A	��p����
�I�pcǏ�YO�	rv�'@�=����5��[��&��!�rm�p	�4,��|�2~�g��Iq n��V��&��]S���pf�*h����x.Fu�Ƅ�`p��p�#]��P/V`
�ǉN83�5����`9=5��4oݚ;u����{Y�Ńq]��MMMOOK��2\KJ8̰���-��/`]Rm���ٵwײpٛ��t��-D��/@���Xik�+�df6q�iun-�/�^���PtXr�F]�7�lO�HV2g'YBlI��h!�9�U���'�hS�|d���}�^����Ԝ�d�Kb-.�����G���jfI0S^����(��̠K��z�s'Y��kV��s����+(��@[Q(P|@=fb!���$W8oLw�L��06K���:)�/j�z�Чӆ��-@(mE~�mj5�-�`=�m����C��5$@�fJ"��BQ|'��:Cz:)����:4�k%���.U�ct��*����ȁ��ų����x����Z&�Ř`sA���Gy��'������y��_��O�����X��+˪i�D�%�YI���;�`�V�~�:%';8�޽��ի�D�+�
�^ܞnE!��9+�q��R�)�:+Y��5�ƶ2�m��]8���m|��'�ƪ�D�Z�}������5�~:���"E�@�h���(j�u����K����#���9��;*��� ���n������S�M�v������ذ�8�T�ȶL�� �2ق-<tm@KMF!�H@+�Jk7��JYA(ݷ��qT�V������[�N}嫣c���˖g�\[8�?�d�(
��!%D�)5lz1�9��J�0�b3v\+m�\�����/�!^`
'E�JTc[�#����f���dr����Wo�[��J�2���b.���6�;���7�_�vynnnccmcC���w��G�����l�^ �BQ ���R9ʶB������5�(cE�ga"� �
�8W4Bv��MyY�b�:��)}���aܭьC�W��b���b,#G���]�gX���˲�Up*2�.� j��#�2m(IeE�[�*�)�Ч���W��!��,�EyK�k���e�v�Э� �^^�T����Y�H��vZݔ�}��.�U Ku����Cɕ�嚮o2��Q�B�U@�Fl?(�9#n��陉Ke�F�z[�¹\�6�j����IZ7s�CТ�V�A�<�a	A��S˴�FO���73�Y��k��� X��	%�3����,c��VG鞭� j�KW�&cR�'O���ז��Ue�<♭N�
��С��q�W�\��YsBeIӜ���G��^�)�y#h�=����,� S6k$h���I�E���ޣ:��-�F�Wp�8��Lv�4+������sqq���g��g?�ka�iN1��74 �?�Z�-��9��c�/^��g�P�-:FLfm���}b�����MR�D	`*�.}��[��#a�nhK�;,'f�a�t*&c�����Ҁ��$�D졠e���U���y�̩W_9�?������Vy�PmP8�L#��y���N(k8��_�N'�7����[�~�A,./T?t�~	u�����#��ڍ�� ��c���:���p���䌗�]�p�}hhx9o�-Ho�T��o`|z���Z���5�Gƈ]�v��du_��� (J~�X0)���q��{��<�r.m��M�ް 8����8Fem�)^�l
����uj\��0ąl
vx� $эV�Ȉ�b&-݉0��V���%[=V<r�<k�P��a�4����!H�L*=:<ric����T���@��El�Z�j�c^��r�~O'a��:P�B.���3Y���Oe��[�T`���!ځ瘝D�3ɘ-�9��(�;Ngo�Jqzs���hU39\�l�/*��m?�ͤb"�߳�.G<�I�������x�.�IF��:��,g:,�I�#��_�"cz$�+��ZF�Gpj�h"jƫ��=�T�ciW��K(��o~��O�ď}���6�ױ;~�W~塇�����2i3;60dс]{~�?�R�=p��C~�7덳o�;�� 	��l6'=�:���� y^?��W�op-:�!�)�.��N�',� �bD�}�!��zDt��4�@�
�n��-��mҽ��_���ڤw�,��:;;{������/�|��-
H_�`2�aB��� A��j�4�"��8��6��F��Z�e"'0�L��7��(nCP@F�ĉ������1�G��{�mF�|A��cX2�������Z��0� ��F-S��诮.y�>�Vb�q1�}�⛥�p�1��_4w���ԏ<���ѝN�P-W�}�Vv�Ό�	iHy����&�@I0̻80*�1�����f���n7Z~��^�c����v���N������r���[���^^7�g��l���j)kG����f�V�N@A�K��/^����۝ڡ{f&GM�3C���~��9wrTU��oM�����M,5[Hka��V�ͻA4j�F�	���w�v3�i4u|C1qÔ���F
���-�]�j����J��Όćq�q7ΫE��6��jZD���Z�/5�vR�<��kh>������8�c;A0���Fi��X���`E�"�T�r� ���0�������ǽ�>��Hs�_׭���5*�@r]���]��f��8�z��d�#w2��}}}��s��j�[�9`_T]��4$fa��0??�~��a�	�?���d�XH0�ɌL,��{J1�h�#m�U�RV9�	M���7�pjjJ���j��ΰ�GՋ��t��ˇh3A�B�B�޼y�$ox���,A�����3m�(�� �|��"vb&�kh�2���7	��'ONOO㄰�/�|��Ϫr�A�P{F�;g��_�n��W_%�Ѥ���_<K�P�N�L*ZN��i
Z���K�4���3I�t���{��X��$2��Y&���ȥh�Ⱦt���	�����^txԀ�]�,�9:>&�Tի��N��/B�`,�Aς	�ӶM�/�ϵ3)r���K�ӳǎz-��a9|�@6��C@.ktlh��27��G��ځ����_x�+�c;w�\��^mm��<x����ܥR�obvP���/�P�#Cß��'��~���5�
(�'�it\E�q�u�u��pf�t*����*�f[%�	�>����P���� �6�A(�y���b�R�Yo5��\1�a��򋯟;�k�.������7�v��h{�2Cer��fA�0�@l��eK�Mf�
1���Zx�3��C�m2��vku�We�[f#��U�Rj���nq�)m�S|i�}�1��I�w�*19��^nXz(��M_��T���2���(4�
�vY�F���YD�e�lm�Aw�fn �$�A�n'%#��V )�$�X$�7N&�� �M�_29��W�b-�7<;��Κ�[�q�f�g�&#�&W�^�җ���.]������oa�ܘ��I��>
��)�<>��������/�O��#?�#'O>������'r�ԩ�qlI/���_z饵��¢�(Cʑ��ܹs��DL�$@���R��3��И����u=2����Bu�o�ԵoIZ�N2׭�򹄠1�9B�I��6d߿��.�b1sҦ�J�LP�s�7`;�u�f>���}�c?�f
���z���}��P_� +)��*I}�2X��b,��ʺ߮�q1:f�
����e-�lZ�Ξ��S����+7_}����`Xm�p��(��7�5[�BN1w,��zR��`'������Q-�O����@���?,.}9Z�A�@�Ǚ�<w�[�L��X��7ʕ���啕�z��I;�|�.Rn��/j��w��NȌ
C�<l��766	S(����@ȐČ�D̺(0�4.�C�ބ�F�R⠎��Fʓ��nڱ3i����ͦ2�N��ENV�'7�4e����9#B�s����Q�k=�D3��3&��m�O��gu�o�ԝ���#��6�EtL� 鳼S��$G������-�+�yV�t�/"��� �==�#�R��m1!D1����zGTr4�^C��P�'��R�7�l��~����/�$\Wg���	m_�h�OXNЅ8	�:�b�X�d�f�0�^��jx���KC#���V�ז`�5��z���ɋtR��pu)�P�A�,1����r,�b<���!�3o�V�1N��5T	>#T����q?4 H�v��1��q�֡#��G�f3ӌ'��Y�����@�*}�333Pc����O�����ݫ�B�����O{c�\�v�߬��U��IE%�I��l
1{���Ì�é�i��)��āLr�-�&�w�{ 
%�c�xXr�qB�ˑ�����X|��Yj�KG�B�}�b��Y~�VY��x���a�|�/R��P�:j�݉Ma�؆ݎ�5�I��3׻x���_~vD�I��x���8v�H����vys���\��jU��VnݺU�l�yq�����v�g�uP�*����F~�V��%�C�Җ��!E��9=5���Y*�MC ��Ͽ�g�gq9U�/QG�؝^�%[�T|!b<-7m(�* {l���j���a����O��Wo\߳g����󅋗~�S�u�������en��7z<F��$w�����0C� �̊!���yinnU����� ��2�E~�U�����6jώu�Gv:���l�%c "OLC7<%�$�g%	=2��s�X ��}\����#�L�+��rǢ����1ۖI�R��M�5�@��9�����t����w|�H���O:qHFG�Y��p+~�.R،�����u����|X���P�j%�-�eԥj��3O���_;�
���|���ٳ�˫�������縟���?��3��?���ׯ<��S?�S������?�������ׅ�Pu��$�0T�k���-!fggg���X�&�c�O#�C�%[:
��,b�-��O��q0{x2`p�A`�=�mX��-AD�
H{܈��?�7|�_J!�u�[���F�Û-��!tP��I~[��_�ǒuw�^{�+/��L<����3���o��<�R��e<��``��?��i���~�����7_y1e��*�����w�H�k�A>�q\%S쳭̙�W����}��Vh�Nfs+�%7[�eGTO�2Q���f66V`�Y����k������!a�H|,�T�")��w���S�n��iHr�������E��v�ǃm٪�������^���Ց���$�p]����FG�R��kRF��,,�_�/�����R�4If��̣��q��2LQ���n��p���C;�ۊ�а�l�nm��r��)�4�$��u�:ίQ�ً
�KL���g��Z�E:K�*Ĺ-J�����F�TЧ���hv�=�$�j���P}K%������Tm��d�]S' ��/�%�����R� {�%݊q~�@#2�%T���R���EE�`�h}���CB�onHzv���P��ٌ�D�V�I���^q��5� &�օ���E�ԡ��t�>|���j�*V;�F��^B�C�1��µ�v[�t]*�Y�4�.�I5F�L�n�B:>����%O�yp��@쇳����:t��~�:4.>d�h���`Q����}��8�9~4<\�2ˡ^�dMLL�T�a�&ƣ�f���XVn ���T��\Z��?n�̙3dgn�3���N $pK�(��a�]�[R/���K�`y�-�$1G����%�æ�
h�� F�uFW����~��Q���*�i�4��Fȱ��0�D�ӝ��,\�M�j?*�*��k*k�kjaXB,R�Ӛh]*nn���7�(λ��S�.�a�Sn)����H��M�;�ʫ�|�Ï=919���z���l>Չڝ���Q2���Aqf�[���ۻsG��@��Z��R�Xycs`�pb�T�[ZZ�q�X�=J�?��?���k�pl5�&�ك*h�#�=���3�^�t�ȑ#X�Ђ��BE�$SFo������VE_)�һٳ���؀��ĥ�v:���K��ŋ��;v�߳���9Z���lK�l$E��@�$n�..�O=����bU���ϓ7�(�*�l���¡W��ի��lZ�Tl��/Uk�*i��;%O��-}� �i1��!0�������\ʭ-��=�X��5O��ڛg) v���5X|O��Y�5������@6]�V^*.iJ*�����ÃC�b�Ѷ��ᴛ���߸I]Z�I�!D�w�[U��ؓ�a���b�M78�����@��
a�ܪ�+kX�}�~��&ӦT�*N���m�޽��]�%$.W���/����ӿ����?�?p����~�/>�ϔWn3 �S��$�$�e.1>�p�{�b�!��� ��qOA��O����U�/bG`H!jH�I-I�@G=Z��7<�O� 7����]�v�s�=����:��J�~���e�fl��@�*g�	�^il#�^��|�n-o�������k��@��ơ����Aq�ϮK��7��P�����ڭO<z����O�N�a'B˄���c�!�.8��d�5���[������鬪:ʘ.�O��d�-.�D�`>۞��t~�GMI�k9$5�˃%G�CL��6j�s��`�T�����e��F1�K�ylOB�M �|.I�j7Z��?�������~~����gϾ����zuld
k�R)s��卡љ�3"�܉Ө �Ԅѽg
5$��	c�NQd4��������҈j�e(ǌr(:[a��I���nz���o`(���m,��e߾��!����6��	��7���f�~k_3]�o����TF��'IO��4�#��[�����B�@M���\X���^���2T�թ�8X�Bi�=y�	<����j��_�R�jU�x��jIκ�v�Q����(HG�t�u�H�<�BB�I����uE�+��� �{bnn�:�` r�\�0}�I�Kh+*'�	���W��C��!����(3dD P�DK�-AIF�D�v<����,�a���c�cߚ��;��c�E�!��ȱ��}upfX3<^��=݅0��8�4���癴��A�㴯������q��q?,�ƙ�Ņ��V�A�*�He�MK@��1"M�a�z�1Ŏ+�h0���1q���7\x��pW��ӰHp����< ���Li�A<,�ܨ��J���:��p)�[>�[����T���P*�����¼��MCV� �vh][Y�"0"�t��T}l$e�خ�]�����_�R����=06ܿ��RnoZ�|���m�n,/�.��X�Q*�!C�oEr�X8jk����8�#��ʕ+|$�pwڧΜv �l�xk�R�
�D@�V�La�fy����|�U��t&m�v�Z}��Ӱrػ��T�F�I����ʲZ�d��t6_^�̩�ܹsv����ۓ?LS�xcik
{]�HT�F\!����@��������z�Z�d�X�X�4���b&V�,���$vr�,6D�mI�4�eLC�t�#��Հ~��0����1=5Dz�2ccc�Y� c��v1V	@��s�A�=��#�C���l���\����#�:�m�Z�f�2_;��"��0܄�8-krD-zˁ����-P�<U�B�li���!g�M�T�$ؠ7�t�̑�0R4�ceksǎ�̮=���ݡd���W��)[�V׀�=33#Eŭ����~���'~�_��/�/����<n�7~�eT<'����8-���'OB�ݼyw��\Mh��~�+����hXQyK�R-:�P��a9�-����ܮ$�r/� �G>��̩S��`E���Bߺp��x�n8����!S��N�hT��p�ݢ��F]e96[����}w��EU.�@��<�񃎔 �]�8M�kŇ	:�LIU{)�u�aBg�Z�\V1��O���9�[����tS�J�Z�Ìc{9�ؖ��6�p&�V��ք+��"�(��'՛A��%������]t�P�[�� ��+e$�E��T&�����EbJ̲�H���,��g$�I��ƺ{��ϋ��:W��-��FU�ݨ,V�믝}���/_�816P,v���å��
#C��+�qj�%p��@���J9�0��-��c	�`P:��ь���e�_m�-�t-�]W�z�>��U�Yǖ�}�3��*�eĊ;�'h�^�P :@ſe�K1Oȓq�A�T@H�+z]���Ȍe$e��K�c�
A9�z�+�ɥ]�-�r��*�L孱�oB��£w��:��nb�\ϚwL�
eR�H�┛Jg`$w{������lXu�(~.,��W�6��D�ܹ�Ek�I��/�|m�p��x��,֍2x0�ih\��?�2T$A��X�F����P�X�To8Z��7�`�6�yY�˓��ɮ�ݤ؞�ҌҌ��}�
��۰��a4f�Ӝ�,.�&�Ov��	�?a�r��5�-����.�F@
;1�؆��Lmv0冖
���=��9,�I�P���Ӻ�ތ���Y���,�rP�8�/���o��L�\(~zp���h��cj��g���ø~���ԙ���c�I,T�Ė֕n\�k3t�ϋ��"�A� SR���F�=뮵\�l���%�;���#���67ױ_�)`����C�z�" ̦����N3)��c9�"%�8�-4ۭ l�N|��]���cC#�\�5φ\.����_���������`&��o��V��HꓤK�a��r̤s�iܸ9�Q)C��)�	|�}���˫+�B�U�)S�4���qf��J�|�ݶ3��H�eM�'^B{um��u"&��1���q��pox�U����}{'29߈�A�3�L6=4з���n�^?}��hB r���f2)No�n��z�U�)�s�� w+��0X�RJ4����ѧ����yr����:`	�V�z}��ٳ��[�䲑�sᄱ�3��\�������#��9���q!J'b�˗/_�t	7C� !C�DS�'��`$aY�D�S�B��(�(���ۮ��q�!���;-�j�B:�~T��&�ݐ�T콞c2�*}J���2�&~"������$f���h}CG��=)d��e�"�(�ź�K��nk#q�!l����o��������?Ď 9|��=�j[������V������>�;��F'Ƌ����|�S�z���{��F�N�Fh�O|������r���¥?���؏���ӧ��~����P݋��p��� �1�P�aQ��̙3\�(J0\�Tr$�м�F��;�p�-9�:`B��p��QL�K/���n�違���q��6�RB�7j�@:�2-�0�AT82��p�Os�X�2'�X��F��/��F+��cޱ!l3p ~h��?H� 6`��F�#�G�[�N��Dn��!2���,̎I:�Vc�hX�M��ז�h� ���J-�B5�҆@V�Xd��ʤ�9oϾ}��Q3t�s��X�h$����}j\��#�&5�ȵ��#�\��\K2*�#8ʸ�!����Rd�4�W�W��91���:�t���3��_�_�Yݪ3�F�v���azGb�xUg�K����R!m�n6}!���j�;;���7 �B�SL��e+��Ro0�i�JaY�FG��|�@9���4󥉣��[=�^kZ0��}Z��Q����.66g�͚��{���F�.h���*a�����ğ,�jB��2����:���b$�.�g�i�)|�m�vdݨ�[��br��~*mg�pF �,)뀬�����liDq�`�.B3{��Nl��eu6�v�:r����|�#�����3�?�7r���kU����T�j0�0,�vK5ś��v9������K��]�8Wft?����I��lX�l�F ���?P�S�0��I"W`�9��V\�T����!>��V)��ؙs�L6�VC��d�$�qb)3�#W��C��z�v$���>��EK
��ܯ��ڭ[�4iUt�%m2]W@�@��;ر����8���ŒԫJ��M��	B"���5XՔz�
7CS�����^�I��E�	L"�>�X^��L&��FLI��?1����i�	s��g��1њYKw@J����60����W�	ei�p��b�)<); q��ED<�(�&�)ݺ����\�#}C}�}�|F�GťRAu�I6��*�J99UG��H8��|
�x�:�A�����]��r���\u}5�W�.5��w}ϓ'~�ƭ�?��Og�Xr��S��Z�Cc�Ι\��������6$0M �!�G�0>e�8��R���Z��I�Xܳ{���2PF������&���e��wS�\�Pٳ5���E��3
a=� ?��Pv�-���D\�~S m��f�;��r)/h7���;��C��͹�b�$
JrFs�s*�iT+���mok�����׷��-㩩��Bؠ(º�z=wbR|��>���s/ݸz(���ow�0�iA�X�b�u��jvW�ѭ���&�&��p�(�߁0�(4l�ՐE.#n:�4�� X�/���a�ܒ���H�y�:���@��v��JY<�f��@H�k{}T���9q�D �B�Ԏ�d�#B8 сs�r�41v
�Ɩ-�/\�@��$+�N�ҕ!T�{sf�azL(K�yl5���b<:6��?��3�b`�>�����36193�s|tr�/��/1t�@_��p~��`	h�7	������_z���#�q�;v��/��#�<r���Z]�1�X��w�:U��p*|�[Nay�������_�"��XT��x&B�v�0 �k�.<2P�W���7��,m��(h[ٞ�'��̈{����[�o�H�����2����"lӋ,l1�J���9��Pqh0�/���Pi�v�R�386����q�L6e۪]ǦQ�
!�ϩ�uǓ�7#��y�D|@V4290�T뭍�r��q�v��=�3?�ԇ=VkU
}�R�X�VW��vaj����Ėo�����B���0�C$��f���L.Yn��'�����r\/�B	�b� ���!5��!�8�J3�t������щ��]/�j�����Q���t�k�V0{������j��,�'����F'g�����+R�7��k �j�2:<C���|�0�^ņ*<�
���d���}
)�ϕr�����۷GoLL끐ʷd���:�BJ-�b�v�t��P:��H<Q:���byz|�?��{W�@�����c�*Q�Λ���
�l��ŝNK�D%�uK�\[4h�9�(k 7��;>l`��� 5!��l�������
�{I��f�:�G��d���eC�g]'#܅�!��r/�u �ڵ����K���sC9�a[����i���S����#O��<��O��O~���#N�-���<��}��o������|�ى�T�KG�VϯBU�X���&�/�|6eaX�+XB�#����V:+�Ҍ�bf9I�$�餯^�ϴrZä(%+k�#�f�CO������:�!x��J���t?D:#{n�4�M2k�#ɮ5�n���T3l�3L(� ,�d��?��2�F��
**��ٳ:��Ňt���gf�E�{�9x��ɼ#]��!��7ՋU��Hc$R�Ȋ�*�=�Љ �-Axi�`V�X�/���0g�D5\���C�=v�b�X�|�A3���Ċ�h#�y>,��i	c��Gy6������pff�i�c�e��Z�v����l�F�J��Mft��sά��+)�tJ
BK4U��Q�ry3;}������P	 g$�,|>.y(��%�K��v��;t�X`��Z�L��Ra(g�����t���Џ�8hv��Ï}�򅋫�_r�xQ����vK�Z+n�es{���M�-�ԚYope�k��nEc��s���,�I�73�b_	���\A�%;~���g;]UY�oTdf2�F݇�L��j��;w��|1�����_-����+�L� Tշ�LbI��(MhF��O<!����}��-,,� �tLMM��_|�����ȑc?��?�я~T�I��~���B�x����K�\:w�\:G&Ɏk�C���W��z���S= ;J$9��
��Y� $����'���$l�:000)ς�wsn�S�������C�aйnij�`l"��^��(C�w�M� �+]6*�l&�:�Tꍦm�����'F&�o߾��	Q����+�� ȶ�N������'?��t��1 ���~����l!@!��?M4J	���bRpK�8!"�耴=� a�
���4�NFGG��o����\�P����?�3?�wߞZ�Q)o�?�h�Ν'O�$N�5���0b^:���[�2V�W������B����� ��i�s�����g?�Y�!�0��h0��������M��!E
}=����R#q��SSd��=����pP�EՏq t|��1�_��W)Z�"�>M6�z�,[N�ݚ�����U����}�{�mwZk��I�v��ͥb����mA{��b�3�.��2�7� Pʑ�,C.ds^h~��l�>�D�4f��l���#�M91�l����>~�}�چlL��j�i�̍"	r���ؔ)ے|?f���rJ<[z˴�Ɂ����\�ެf�'�L�ĔV�[|�∌�w�'U$¶:�;ܦ0�@��:%�cK�a`�uS��n�ۛ�j���>�F{�ܸ�x���O���gfv�_�b�O��ǋ��Qz���п����F��̬���dڳr��-�X"Rj��ԓ�9e��˛�L>��h4k�GD�\٪wA�.�B�m͖/d�F�0�����[�5���Z�T�܊���j��u7���vտ-0C�(H������z�X*�8��/�
~ʫ��H3�<�b.�1�n._L�ؽ�q �C1o
���/4Z���?�S���o6�>.� �2~��`�T�//�;N6;d9��F���<�݊S�?s�$�u�	>�^��U]�C7<A#4 	�!GiHJ��rW�gC�(��~Q3�bC#E����Eh�\����H� A���F{����+}>�߹_��D7 �&D���fUV�{�]s����@�B;�����s�Ν9~���y�F�XU7��(����lG�B����3��x< �$ܛ�*�OFK��g?����Ooް���������������/��?��*����k57�T�4Hv�s��t�P�:
6S���"~WFn��0ܯ@0��&�a* %U�)�Q ��Lc���+L�a�&m&ڲ�U�i"&�Sћ�,)HL�b�S=B�C�2)nqq�-;����FT&�	�DǸ����(��3#3�� ���/���<{�����ʤv���	JS��[�8qj���1�g��mO��rF���m=Y�Î�x��B�sB|������;x� f�e��H��CH
�����E�;燾O&���.�9s�W^!�����-0�:dǿb��yf��(���mM�G<���g������]#3tL�\�to<3m��&,7.�� RM�{�`��t��@#]94e�"�S�4g ���W#g�P�+*�pvr:Je�a��3���A
~03>Y_ZJ�1>gy-��ꑦ�Q��J.M�pޢ�c���r�Vod�={r��]���]��R���̉U_��J����䥫Wϼq�J+�ů�vdaa^�B���s��y&���H:&���	���W������~�\��?s:�ג��_�T�(]^\є_"����y�R']!���dyA��l�lc| c�7��.uBm�พ�V����D�L�::�ƽ�Z�Q_��2RYi�QW�o2�@[��v̶e�0�!qL���/���ܒH	�����G����W����ߥ����)�wK5a3'� �����i����=��7�1�935Q��n�:{�R�����(.: ?0�DP�I(���
0����Kc�7�r�ݻ����	�MB8;[(��С�q�Ȼ��v��ú0����U�'�����*A$����>}��G>+V+l�����y�3�Պg�+_��'?�IiR��3xd]���<g#YS)�}�1���xS5t����,��Nse�R�Z��7���v��F��P��+�"+Fj��/_��w������m�H�(�à9��
}�o������x�P)8��B`�R�+e���`�^{�5</���� �:�Ѿ�꫔�0�:�OҀ���� �jj��b�(6�6�M����z�A���鼆�{GSY�_u��'߲٫~S����΅�B!��S�ڵ(z�駡8���O'x���v��h�p?�y���W Q%ġ�l˰�r�]�,����9�b��{]�0������y׭�	���>i��R�@&�Q�g�)2u�<Q����G,N>�0a⹁W*�n�����-q
0AJi�m��@�w�Y&K<�=�?�幪?����f�LG�0&��{qn�رck�U5	�Q�XU-��:���I3lI23?�GF*�
;�.,�8�CI�vJ,QX/����T_Z��{pӆ�f/]i�8IkݮGeIh�	��ŋ�%���������(��d�K�q��Gbx,���&L��oڮ�f+���j�k$���E/8Z(Ƨ���G�4%@*�{TT��� �Ųq�rŅ.��Z �ʾD�Z�����ʖ��5k'j�ċ%a؃�5Z�(�ڦ�� ��~& Lv���@?b	$i��i �P�
��Q��M��R.L������v���e�����l�Z�ÀF2�\S�PS��.lVH����������Y�{%G���������=[��ٲ��u�O�pj�΢��KT�<gn'w��ޘ�UB$�~ڧ��,玻n�ҿ����k���u�J'�N=��K��o���-��}�>��k'a���\|d�P�N,hֱ�	���U�0��� �6../,/	�.*fj�at�N��ғ9T�{�4o�pj���B�IOme\��M�X��n�s��I�{:�����(�w�r(���VR|3�3��Y7���Lq�9�b�ѿŗ��7(O1 L!�c鼦�cm�ѣG�HFԋ�SZ�0��	6DYlL�-� ��)"܄����6b>���'Z6�/_f�;K����,`TsF�F���St����&�031~rg��Y�\�A��;�ON*f�0`�w�1L>!
e98�.f�=�y��ݻ9�ddLRz�(��W�xK<s��y (L&G'r���i�s D����MEq�u3��lx</ߺ}��J|��d�mbсC+L''`p{����0��v`�J�i��:r���ľ�Y��]R9]��Q��:�;�Bi�V.%����Ԇ���A�*K~Y g׵?�
��\�7��$WpU�#�X��|��ϢM >�L��2#�_<��X�-,G�ͳ�^"b��\rk-��n�9����={Z�Gߠ�%�NϏ�Dp�m�#9�Ʊ{V��`���/	Ŏv%��ٍ?������?^^X�"�����%�#FGy*����>����w�<26��Qz
�
P��Р�ǆ���K?�Tk�$�gw[h-U����'��O���'�w�*Af�'�w1?6*[!��o����ꯎ�O� �+��F���sj���?�O�4z�����g
�%]>'�r�-�8`�N�8[���o���?���Y�����B,@Y���ӱ��4��i)u���� ��4��q�_o�l�K�N�nm�	A���٭;vL؎u�Xki�-r�Ա��m�p�1��=�}@��~����~�.���N�y���B��k�5x��+��yq��@��S�W��g���''�q�x��_�Rhk�}�I�n�9ì��$7o	��2Y���}R?��_�߼�iwם���=��o\�t��&��y�ůs�k��Á7ΕdD�կ�V]HD�ؖ�v�-�bK�f��ssgO�޼�V���Gz+��~�����ILb���"׎�i��A��H٧ce����:���-�����åb�{a�S�a�65��f��6��o6r3T�Nn�4HG���l�.=��G�y���7��yC����3n�o�4cOŭ�T�6;a��麥
3�1���/=vBx�9�w�qǁ�XR�a6��&0�s�W_|�����_�P�T������
�_�Fem:4Hu�;�b��^Գ=�mU%�)��b%�5ǧ��S�8>��<ƆV�<q+G�T�]��4:Q/5������eSeŬ5멕��T!��v�����$��[ �SĿ����Ɇ
��,�
� I�uq�%@����)�S����K���	 ��9(�05�0N�#-ߍדn�n@�x��c���u<_��*���zQyd,��+�6�0˃0-�I�7T�ԉC��]-�##��?t����˫˰-�J��0�gI��!�w42	�r�9��	 ��}��o��M��/�|�/:�Y5_����O�/�?��-{�:~�J�k� �%!C���b\J�BQ���s�gL�U�b��9(�a��6Xy�u���{b<�J��:X[�Z��L�"0��H�A�ɲز�7of/<�4=7`{r�����i:�d'����LT#�ќK�,+�8*��O�>�_I�pY�R0a���`�͋���8	nMLHh���n_��V>]�4�Y���,���`+�,�_a�1�ԯ�Ǐ��	�<��ӌ��sI�$��|R���h�S�A�pW�J7Ⲹ;�c� ;V���p���`�ur'�*ҍ��u�,l,(Q���J��Y�Yk�?\
�~���[1�&d׮]�l��	x�%���6n܈�� /�la�ӎZ,rQ��Ew��4H�����\L[�P*e��:�Zy���8�:�ȕe���|+J�N/i��W�|��r ��,�L�Y����];V�����
� 8ۓ�i��V�pp� I;��tƐ��Ҋ�o:��dϪ��M�R�?}K�ϋ�	JBT�����u��-�ߡ �"��!��Wr��,�ܖ4�E`	��/�rY��_�Eͦ�d(8�a��u{r�lޑ���ښ�/�e�V�=(��~��c�|��4TcM�^��)�H�q�+W.c5�����_y��s����Ɒe�S�M�*R�C�z��^I����JE�r�^������fo����8�S˕bܓN���b#����S�Ơ��Y_� &�e˖-�2$NƏ���C2F���Q���vo4d>uF�5�g�еlnl��09�Q��({��J :��lN�[���K�j��G�]���K��\�6�;�j\���p���0�r�]JI���Ũ+�S3W�VV֗�n�|�-��V���!O�Bh��ޮX���@{�~�w~��}��7�t�����^z����f}}l|d�T����$B�P���rn��y�U���g���믿�9]�����d;8
�P�R����;e$;�j�Ja���¦o�O�O}Q�t�x\�y�QQ>s�B�B�cJ_}�UHcJ�oD5�-�.��ڴo�:�=���S���Lr�M��=\*��Ա]#�}��?���t����*QVf32�6�'�yt�_L�y�����Y�f���lu�WĶ���sԮ�,7:������#�><�����a�N�M����L�2����1[d�m���Ay�C ��5�jJ�3�D�I��z�#/�����'(��JᢷN�s��Um7;Z�f�w<N�l�qak�x�ܹ?��?޳c��Ԭ[�A���En�ū����r��{��-VʳS���s���pb��rE��Ä�&j���c����ӛ�͒,����U��,�f^o�C��7֮TGg�9�J_��b�_�H�_jS� �6�(�t��+�9�H��m׷�G�t�'m�lHêJ���w�Քh�[������|�D� �;J���I��9���a�n�E���,5�kxN �_��b'��m�'h�B����-��)�Fj�Tv���ŀT]6��-�26�	���mb7´v�4J���5RJ��<YX����D�+�YJj�����Y�� v%�$)δl�*��Zw����_���G�=�5��{�y�]w�b�^ki�����3e	�/H���[lǬ��T��{�}����Au���N/�7s3g�ކV�0�n���5�E��u�NÉ[�խ�^�v�q�2Ic��0~�y�E%&������Nj/�6��L��G��2�Eɺ��V�s`���é,�j���<,P�B�`�B��tU.wF����;�JfK�Ű�n"I�7.N�]���eƑ��I� �`��5��#E��P/�-����%��0]�3��r�u���,�!G6a_,�"��Z��U0l��3G��$����h/��D;ԡ���><,Ca��̙3�o��2�֭p��R�|!7��b鈙.���r
�T�4=��a�-V@��	d�>��ꍆ�Ru��]B-�^au�	Y,�-��[k��i�pC�$3�Y�ދW۝�$�5���q�~Qq�tY�����x��2VM��4��G�4�U�TNj��0�H�g7>T�=ge���Hm���z�x�P���Dr{O�,����^���X.q?��-�9P���� 7a�RU��}��B����}�<�Գ0��8ĳ��اQ�d`b$&�/��/�x�	`6�<��ݻw3�/�<�� v4��s�����۱�l!|ojB6<e�p�K^��$�������-�&�j5���26T��p�`7c��^?�����#���TI�ə_^Y��/�����Y$�m��i�����' ��~�����-�i4���!>'A%N�S��F6?��
�GR��Ts!�F`BBJ��p\���}L闿��|�+���g�2DY�  Q�p�ΰ!����!�8}��S�$}6P�umu����X��P�E����_�Xn�ܵ�����nv��Q�G����'�&�&(�]i�֭'N��|���v�!'N+5r)W3�j�F-� Ieh��t�M@A������-Hî	oH�y�l/Fx��JF��M���=�4��\�Nu�D57B���0/�\�p*�[m����r8F�� �|���'N<����g�{���I��Å�z�oWC�v3�s͎E-�$d�z�D��$�?��ҹ˫�����w�X�c�e�I^J�哐��q��V`s\;��S>��Z��I)Yƴ�˗�a>��v������s��(�).�6���e�&,SdC-@�Ԙ�S"����V�3���n�gϾ˗���ֹc�n9�Ī�_��@ʿ.�S���f5�i�C=L�Q��W�O�O����O<����F��tLUD��tS���n�t�+O��:����_��'>V���9E������f ��`Ҙ�fi��վi�~��!n;1�L�'`sJ�L8�%JV��:w�kޮI�?�G�L	�3��KK>��z��o�% {5�Q���H�l��{�
$0KUy�+�zQ�#����:�8�"ybJ��a;�Vl�a�d=�J4�4��4nw0�^��:���W�Y�!q!�|�, B�%q'TP���,�Q��*�[�]_���\�9���M����T�E�G!�l�+J͸׬U ��D]��nә���@��6ÙҟP���h��\��\��=wo�Mm��^�:����[wM�]|���S��TJz	�&=-��]U�;g�<Ԍ
#��^�����J�Q"����c��=�yAݙ�%�;�.�M�a������	���,mw0vIĬK������
]]�Β$�L\W��C?A�]�|�tt��8��F�L�M��4�ݥt�S�Ҷ֔�zr4K��e	u�D&q1�C�H�@���p;�y͜{>��('s7�^GZ��c���7��k����X�%�՞npD{T�]"��C�>`*���g��ywM+��<o�[^^�l�n#ؠ� M#~:p��%�"4b0�%�$���2���Ǉ����a�0�&&�pj�wF�����4�Kɐe��,�u�YN2�J�դ������F��h���F�hF��J®ז�sn;)4����j��@�J�V���rI��FSlz��1a�.*�!7T�a�ɵN/��d��=|�Ra�nO&�Ç�u�]��K��N���j�Y��L����V��%�=_:�E��6��Z����j ��������46:B�i[椸eێ���_:p`F��ɓI2/d�ʰ��mi��Ѕ�*�=z��#��P�txcr�j�'^|��|��;0�����̓m��Ylv��X:�J����ɓє�w[�Q�4ZY	�d.��G�"��rkv��_�/�]��V;U}|=V}aaW�R�D"��7+��i��~;�~��wR����m���{�i"U:�<��5h�b���ƀZ�ӓ�N4�5/ec�<��:�|iv��":}(
h���Q��5̏Lj��AC���p�H���ϔ8p�RsY�;��[v�w��KG^y�����vM��r1H���+�K�vf�,���sg��k�c#����B�i���2�"�*�"}O0ٙ��:x������ꫯ2�̕�S�-�1x�Y L=�P1u,�dj%3�YTIw�0����|��5�%�L��X�?�5�0ÛF8���]Vs3��t�`�.��8��N�b�	�XT�E�� �=��h�����Ć�'�Lq�ྒ��!n�x!7�v b$=����m�>u����������Daݸ����hQd�G�+��.��G]�{��g*>.?�rܶ����TE}����A�a3��½	�{��ʂHLi�h����ev�b%�b��k��7b�f"I�?2�fv+Y��
�^�O�� O��ٍ[6LXyRou�D�9y�݊�c)k�ew��ٗ���Z\\~��g��ޮ���o���҉���Ŋ��r����E�G:�_�׊�M�ۜ�#>u={����w�H�o��8��?��l�P���P`Ҟ���l��.F	 e\s�Z��Zot�y�N'�l��N���I2�#��q�=����-�P���Y��\�Z.����"�a?�L�R��c�a7^iB+S��T�k��o��R�:@�r�T
]�XҔ`�d��#�	C�o�뤦p����,mL��Ŧ�0��M�Hydz��m��cQ�٬�F^r�����ZV�`.�f��kt{^h�6��v��7o�x�T*�?�Ĺ7�l,\�(ID��;�� �6���q��~�0E��)2��凱	)Y`�h�2�+ց��������Rw�cd�&,��ä��v7�"nMjh�<!�ڡ���A��T�A2��H(-]���^@�4$ǣO�#ޝ��ԎD)����E�n��y;��G%�+��A�5� ����?�;����c���X��bF<��0Z�21dL@�%5O;�h��W�c�ӗ���d]ÿ|d6W�n b�ˍOb�0Ϭ�cе:�:BG���5��QfF"��ҋ��~������ �#h��I� �m@G8��r��
ȝ�/�P J�O͒��?�R���{���ו�5<&n=3=�45		�pHu��h[�+4�I�*�R�*d�P�����"�����Fs���z�$7�Hm#�t3�a�%7pmU���InK���l�>�j�������;n�����/�|��玟z��#�Ϝz⧏�ٷ�j|tlljjey���
�BE�n�iR.���NP�C
h�x�BPL�tiqa�\>w��g׮]����o�yrj�}�����?u�̓(�w&���=*dc*g,��b �cm��ʯZ��+Ele�w�Վ�Nq0��	KPR�:8�_a7�2"�!�گ�ʮ�y��X\-+Dn��\�!���&&&��N�>�g�fS��N�\����FFP�����X!7���Lz�����\ LZ�f�R.u�%(���T��@>)��v�0�'�ۛQ���_~��7�`YnMTOM����Թ�ڪ�S�����}èe��G�blt;KuKe:�K#O��: �0͸��r�KI�f=��=�q�w��-�Þ{un��_�:FN�����q`���j��޹t��6��؊$�Ǜx|�(r-(��t��x�9f
:JzpX׊7)�X��u�n��	�����1(��d0���:O�5`0H]���3�,��,����]ӥ{Zh�f1�r�US��:|t]P���~+��Ix�@� �������ZB��Q3&� �����B��p�/�*Q���49�g�k���x��iE�{���	��(@i(&�w
%��.%��6����'���Z����b�I�zQu��4�c�z��3b臭~"��o,!��AIeڷ�N��}%e�,7 �a$?�5�U9A���ķ���v�f˻��r��l�GK������+q�yf2e
ǳ�ݙN��n2m�ܸiS�ޛ_>�	I��燂Xh��<�h�����\%
�8����M����#�sa�'���(V�t��.�竓o����*���ܥ�7�� �(�۔|
��b}㨳��8wy��{�0K��mb�
2>�:�zbG�ְ2�V��`��@21`u�F��H-�4}�#��r(&�h$ծX�E��I�n˅\�iT�$�'�N��Ҋ����$6�L6��y�Gy�Q/%(0Z.����S�!M2�m�?r{iؖ�X¹�e۾#M���0�U���붫�bm�(��᠇j�Z��<�*d��֐o c}�c�4�XZ�Vg6l_שּׁ�"{�k8��W��۫W�^����ÙF$�*���oUdj�B��&EMO���ք����c׊U�W�S����9^��K���:K�4����(��)}ZTx�'�2���bo߾�ښ��4�1�����a�9P�r�d7��̰�������������(�Y ���t*,..^�p����L���H��׫i����e�s0����Ll�W����.)�6m�DNht* �MKU�oS/|�99�.)\vM�]�@?��q_|v����q!
D�ru>!Q"�������q�����Ƅ��M	��&J|�����N2dn	�E��""�����Mb"�=RZ�e$�K̈c��Mx|�kK堥}�0��6�t���j<�-*�)!鋥�+Jbn�+ﱈXY<~�T�UF���%ڂA�Fa�M��������@8v�#犧�����Qd6Z�o�|'��Q�Ж�M�8!兆��Á,�L\��wأ�+�<3

1�&Yv�$��y�Y��M�RM�{�G?� �f�X*x>����N��f8�jw�U��Б�"�P)T`�\�x���G��0��x�{>����'�톧�2%����#Q����h{9�C�f��ʅ�*�zwl�m۷ {b�^�p^�wi�����~�S3C�4��k�.�o��D;!}G1T��ץ�K�	w{~��T^�|vz�_���7ߌY=z�(N�*#^rw��{݋�\_�&�����>p�M7�+�?��׾�5.
7�M2%m5V���Fº�V�R�L�����a'��}b� 3H��5�wt_cz
��&5=���L����FewQޗ.$��UO�m	�2���t�B yU��3�<��W_}u��U%եӦV�J�����KK����X�o}�[,�Űtu����{���VS���Z֫�C�(��8UM/ ^06�]�I˄NG�˚�S[��q��)�����`툍�tx1M�1��TN�loI���CQ�A�F5��E����2�Z���aM?&�s��u�a03Ԃ&N��t�:uJS1����N�M-�;bky8�[�[��|
�}F�"��T6힄}R��7f���h1��r��$�xB�W��l�DZÊ4�Z �%�APKIOzmNxd8oP�q�v~�ca��ӫXL�D8�p|�h�m�,�e�Z������Z�)-�i���@h������0��U��uD�B�ʉم!,�z�MC/���)�*$���I�2-4{����a2�8�V���U.W��Z�iPs�\Y)����bn;Ri�j�5h��$�/-6ɉ2R��i�sB0`X���'&�KQH�����!���ӱHo�)B��X���0@��M��fT=�؍�wÆ����4^��*���Vc��=��[���Z�]��f؁v��
��H�V1��R y�8c�^���9� ����&�NbH��QeDv��w��I[�ω���,����J�0�k(�8�m\]k�ʂ�Yib&�:K�R��u[Nn��`�\�qصR��'�v]���:a�M#ò�n�>1:��f�I���
�D��7���M"df�T����ƛ���=T��X�)�Q8p0w�d�F���y��m^�;�ru��Z.�(�y�5�-�[�!>�(BJ��d�0����_6T��+#.�j�v�z�%��I��uO�Q@�P�b��t�C�-mbҶ��{��a��J�BCj�ud�f�>ƤyJaL�?w�%ʭ C@���ے�,5�<{_�2�@3%h���� ����S�I����9sF?;K�``��9Ms�˱Y;�����5���m�VɄF@H����t���tT�<F顩�G⚰�Hb��G�]pG���V�j��4j�]����Vę���{��ر&��yϞ=3�ʄ{�T���ak�j".�R�:0��֭[a���'?�jb�<�?�={��9Q|"vy'��΄��yL�e� t�ڣ<l��h-'�Dg#��Z-w�_ 9�wY�/�ʓ�tGi�g�ej�r#)#��acx���]�r�$�)�j�*���T5*GI~�T�&��N"|�B�#�qŜ������D],6�g6jgض�TpnJ���sWz�o��cssW�-A�gΜ:~�1=v�'>�ɱ�1���1� i/b�x����BF����Je��Bu��'��}Q�bK��&;�0Vl��f�Ĳ�B�0L�@C�V�}n3bx:8Z��z}�X�8�����_�Ezv����l/I�Ű�� �!�0�`{vIj$��~�E�utj�(�1�	�eKRٲtܺ�;p^x��v
��#�.v�uܸ�Ĥ卑+�Tg ��}/��O<�=���P��(H��T�YoH�7���-�!��H������ld2_�D������M���}҂Ci
��E9'�K����d�`�9�aS��;���0�G������x�=���M��l\�p�{��ޥ�ՙ�|[2�1K�s�lX�4��v���~�R���c5�/�4���7�;�LSU�c]>����/C��Q�e>�z���:�����ʅ8�<xd&rkb@�5����� ��q�Ň�~�l��`��Ÿ�4�\��ozS��\
:��3�[{35U�KwP�k�[3yA��:�aӤ�/�8q�y��@�S����4iz�t�	&z�X�s��Pޚ#�R�����+�/_����.]yLl��0T<FZ(�/N�Ze2�r��t�=�!p	wwATb��C�ہ�!:��^!o������Ӌs��'{�+�Q&ɱQ܃��9�u3Cv�>u�D�H�:��6�cd����X�����eD��"B(����2Hf�hF�TQ����S�sG��R��JㄾH'��(\1B��a��*X��0Zb�`�z�fb@yBt����<�|����7�r��sBf���^Ȥ�g�����M0X`��w�q�n0Y��2Ʉ\[�|�2� �����L�D�+��[��7��V Z1�9I�|7@������{�����g>zǞ�3F�A�����,�����6��m�� f��H�<�z�Pe=���J>�nɆ��Z�z��ߩ�;ء�9Z-$�g�vq��k6ąY�&����6>2�P� T��5C�}�ڈMH�-L����!t� V%Q�~V3}wyi!n�`J:Y3�+n.�j���+ކ��$٪�QOЌr{T�c��� H��!3U\Ȓ�'K��,�YPc� �Ҭ���fń�[��j�#�Bea�4��r*���{�I:�'�tWN��v�m�if�F���� :�c�3�㶚��d��a��rm�� ���#�j[�3hjc�U�,�a�R�i��B�W�����0���J*u���*y�����U��е�.Y�6)�I�t)���&���f�d�	�5$x.�*����<V�0������ˢhܳ�݁0��f�$}+� ���4qe�I�9x8�<�5>�a-�K�V��v����pM<�JX�"l�7�c�E��rX��/�KR`�el(B�FZ0��;w�}W�"�#�D�FsN�t,� ���"x|V3c�HtˢU&/�ȃø�n�m 0�F�V0��t4;v�x��ߢ��L{�uQ�VW� GE�T�$uفq(q6,��na��6ώO��/.98�X��`��qh�B'�z>�"�t�iYi��[p��`F�L�shD~!(t{8gr<���}�i��ŕٙ�F�36>�g}B�CŔə\��g�,�m|������W�����Y�Fڷ�3�'Q=O�b����� c�l�˥�r5
0��@W��������Z�d���8�C3��V��%<�QXp���\�4��k��R�]8s��Z{�;nߴq��R���3����_q��������@A<״ڇ9RuO���l�R���=۰|�De�,�/�ݹ���|������^$n/̤�KJ���{q��P��W��4�y����a'\_]y�����b6K��:��w2��4��Ɂ$�|��߇���^ ��_~�]�k��hT�eV�M��o�Tn����C�����e��˿�z�;K�2�z*���u���a�"��&��f�|������?Z]_��qZ�;	����Π����X�p���w? ����������)��.f���<��K�<'��nf̄̍�7Ҵ
T$�htd�j��^���>y���S`Zu�	��o��w������A���=wcb!( �7l�b-Q
����T~Q�s˰�+�ґbaL���?|��W����V��v�ٰh�f.!@��<�4k�3�R]{�xXX�NNƅ E1f�
{ {�#dh�� ��3��;�p�����Ŏ��*��V�4�E�kRw����G���g�#G���}��H\�)@}�TI�҆Q3��h���[hLeg7� ����&�J���@ߺ�[n��&J�
0��+������t��:����ؽ�k�o��K	�tgvIZ*�C����jva>A�T��/�KI3mI�믬wk� ����7�,�0{f�g{qSq��!�b=�5��J�73�Q�	2I��i?�kK�� ,JS�$��A1u
uf*.(�FI���jz�:>U��VN"e_Q��$���˄}2��-����P,}Z�q����C�A�c��NONm�ݔd�������`&1Ez�hR^-KGA��h�x����k��ֲ��K�u����Į�����J�B��ұ��xV��Yr�B���=�� ��	;�(6����ܠ��n�������ڱs3���/�$�����g<H��u�~8����SO�Z��T	����R޷w�Ԇ��{�+�3�5���Vysڨ�{����D���N�qxǁݻ'F� ^�5%In ��K�I���S�i�s",j��]`-�	"�	)ܜ��(�PY���0RyhvWH���F���n�UA��/xQ�G�P�۾8I![�Ȩ��V;F��=q��[�Y�eӼ,�Q�ٍ�v�L{��K绍$�2��2�Tf���
N�rr�Ɩd�#uŹ%D��ѧGȯoaX7ά��
�
I+� �!PzQ,p�=r6$8�H�5m#�k���/B|����	-�#��$��rW�O'��k���H姫�ub�v8���yGL��j�e5�]hT���1W����tȝC�û�M:�������at�1S����$���Ϊ;�v���]�jcb��O�+[��Јx���9�	d�O���x���.]bԋ��D}�8��0���M
���\
Z�v<�N�@��1"�nH\�H��.j��X����m�6�^�>Ą*x��i)f�0 �ŷ�\x��cĹ�yxvF]�W !\�;t�2{��&2�O�[H`��5�w����&�����:+���S�EQkr�(#p%�/��t~&��S�&c?�%�fü���5e�p�(Y�v�O+����f7W�-����=�a���I�b���ĶP����23���q���Z�=9H����05�]�]^smtbtr�L�\ó�S*�N�h_�u#2Ǩ�E9�	���\���b��5���qw̡�e�s�Y���7������+��l���8U��Ӱ�0���� ��}���&�W�za����������.^:t�P�.ϝ={��;;��s�?�y��r���]l	,�3�{yH5�>�F���	B=Y;[U����p�z��4�j��H���l6L)Å��\WѺ$��B��oO>�����|�C���\lHƬ1`�._H��l�$i��N�}�����|�G?�Ѿn����LHGso�,�}�G}�?��?��>����:��[�.�Q�\&��9��
���~���]8��ѝ{w]c�sc����M�� ��lX_[���~v�ԩ8N51��§�J/�p�MJx��b �6,)���gJ)����ϩq\����V�[�7�è�����O��@O�����b� (��F*RNU�)�Jc��3գo�?����>?2:�;�ȼ�豓'O�m��ҢC�\�6�&�d*����&� �| \a`���T�,R��>)?��j5���@�ؙ���{���N�`>}C��M� �el�CLu��R<��c޾};�!d��ӧ!@��
�d}&{ӡɾX��V
���qo>'G�Y`�������_��_֬��=�رc�`t�;wc�m�qd���N513t�~%+Qݑ��.\l��VFG�Gj��%!/��^��z}!�{~��[I�[.V��8.�IɊ֔�qie��M�䘸i�Mi&	+&ՠ�����1ۦg����z��۰�I��>���Y�0p��j�L����pU���]Ǫ��si@�5
 {�,Y^]Y[o*9��l����L���AJg_>@�f*=^=7J���/�<}foP�UJ��&����$oK��u��A���Z{em5rs����φ��-CȜ�$$pd+��ᕊ`�,7��ז-{�?y��!��}������Ϝ5VV���݉��=���P܅~v�>�?�:�xn�b�4u�{��|��鱉�ꨣ$l�菜A H��X{�$��|,��,eAU#h�t����ϲL�1L���Dz���Csw[]EP(�X{�M�]Jk�IQeҸJ�i�FPy|���ji��ܑщ�;v�߷��CФ�W�,�� ��`��B�,��(A�3�H�:�,Uck��0Y`v}+=�ϯ����f���=�Z�ɝpS��I`��� ��E��QM���m�B�B����:��	��\�g�d_�g7�jE��V���:�Ĕ��|��#:/yY]wK�Gs�Pk�Ƹ9ӑt��a�&]PP�9�b��ߵןN&�/GW���^:^;���Â����"�F�!��W���`�t�,D ��������v@�0,����e2=`��o��w߇�_1�#���	��+�XJ��"�!�UlD�����c�y�Ö�����dv�ƫ��4Vxƭ[��[�sq����Zgg|h��\�8�5�2�W��a8T��q���={�Ձa1K�m��Et��p%1	�M�|���ώ�4M,����X���K��T˩�ڲj��k'�ۑ>��VGţ�Z��# ~3Ӱ�H�
,W鵎����yA!���ѓ���T.�߻ojf<��k�*p��ga%���U�>z
�0�MW�R٠�7�	�-X��gܾ}��߹����s��c؁||�pY̭�jN��1���s�����=y��ųg"�݆G�gn���];v{�h�Z���tZ�kuu]|��%�{2#=p�&�b�_�~�wN��^]\8u�d�\���6�llu;���E������������E�ZƼ��)_�!:?�5OO&�PX�2�C���xIE)��'|��ay챟=��3�����������nZL�
�1���h�4�����VG~��'��q����v�X*���t]� �ٻ��{������'����[���(��k��pE�)�|ؽ{���"�N��?��{����c���ت^Ew+��ܱ���qfՐ&1b��C����a!��B2`�&���J�,ͩ:��������%a�j��r1pK���ե��������rv�,ɔ��a�S�U�HΌxDM�,��l��v�B(XZ���� ��׭�p֨n��y $�&��ؓ���9`*?S҃���p�PkkuU��+������H�3+��w��O~�[n���ǂ�A�@B󿳟��X�F���n�	#�t���s�uk:(u=�Q�Q�q��'lj&7�
`�%n��/0�6�����)_���7�.'��HILx9LK��+Q�.��f_o�	+�r#�Z�x覽- �^�:�Jɛ-�~it���n�A�qS7����ը�����Z�v_�*���M3�����4M�\Y��q��C�B��:]�F�ߎ��0��}���ʄ�5�Z�,��]i% ��k����Y:8p��RF���R����?5>����%(�e���]z_:I�F��a��_UD81%s*���ة�3/�T��B �|�Y�M��Vk=�z��`Z��y%0|�yb�#XJx)�4K�,4"�!�s0O�)����mI:[Ҝ�_�r�ȑ#0�J�r�Zó��D0>K�~�s(D(k����6�.�ҟ4[m��,] η�X,S����*˥yVvM�X���ٿE#0�˙�)��i|�����U���c��P�l�W�d���[V25��Њ��������Ώ�^���?�������4Za��2ӳ�'�v�33&��� ��#	����<UТ�3�݅������I��l�1��[�2�
z"[zQ܁�0T_##ɆܗB4����[�����
�k�7��vZ��E��㵙驩�^f;����ݏ�\k�5TG�5�c^�F�Y2�Ȁ)�@� �G
Җ���#�$���d�ݶ�����/���Ⱥ���5"��1,3e�,��LhP*� I��"�=t*>F{ǌ���� ��|LW�*����a��ݻ��c��T=���^��?���zDG�����z��X�Y�DV3��V�S�p7��H����ؒH�8�����x���ܔ��� 2~�4?��Ic�;MID|��c�lB\��1���|_�t��\*N��Q2�*�A�b93� .��b���E�qډX��,��rCH���7�*�u�]+VTZv�����	�� �a�f��$Jwi�{�z��a��B/�_�P��S��=�v����~�ĩ���YJ�T���]M�Y're�ި���9�`׮=@�L2�݆g��$�i��,�={yii��_���s��ǎ�������O?���-\]�3}�c����?0�O=�l��Y��w�����>-���#�vza��~�� B_����⋟������?�}���w�u��N�[d����R�v(i��:,Dl��-�]�r��Ś�z4����յ#��:u���@M��M�v��[��E���ܶy���F��s����h؋u�t?I{@�?\�*Nl�p����<��ѣG�N��]�v)��uܸC�~�W^y��������w���?�)��p��k�e�}����u�܅��!�g�{�����k"K�wZ�(¬�ҍ��v; ��r9����M�n���R�u��b��,��ѽJh��LZ��bOX�1ƨ�}mکj���;K�T��&*��Y�//VFG�,ޱ�,�1�vm����SJ��ђi�ą�6P�!���ߛ��z���ʰ'kMr!S��D�FZjffg��&�-LKn���1`l��ׂm�6������l�v��r�Ry?�gM�������?�-�SL�RJo� `��ŋnl�yH��;�h�@_gv�����C���@:ָ��!o*��P����~'�nDH{L�n��J\
:Bo�%@x��t�t�y��16є�"�'F'�/��[�����̧z���O��҉��^L�(􋒜��!�r/��$�v�����h+r��n><55359�aB*(�)壯�r�ɟ=��O�뫞ođ�M~1��oo�f�OFn�<�B1H �̬�"��7��Yvm�I/��-��~�t���M������) ���LśC���c(�b�͠b0��4Af���#o���45>�)O��������\Y�����n��ܖȄ��9���N�.�R~T�%*�R�s<;�a�T:�V��m{�:�P����d���zP����0�yQ;8׃f�u}�A�w%b��KA��a"D��6i�m8FU�T������ȁ{0�����FPr�����N��KnxE礒��>�_Yմ%�ިd����d����n/�V�f#rc�Q�j^�@��l��R�u��Kz�bW^@[���>2��ԇCd��m}]F�b ��!�^�ګ�U׭�V�i7��Z��)�;&�!�v�:�9/H�"&�Z������t�?��?�LOn����k��
����Xbk
6g��WFl��Kǵ�Ɉ�{��Yj��u5T* ��1,G&��"��Q�ĉ�:,Te�+S�t;yMX�	m(�5�Q�˙3g`Ѳ��?qA�Q��w�W2�b��X��v�+���"�*�ݘ�����X,m��I�����;�<F�AB'��9�R�2b��x��p����Ӧ���ʖŭ�;�"f&��m6,|Xhy�Wh�P�g��QI��Z��W_� o��f����#4f���bT�4�I.�tqe�f����`"
��t��Iގ)p�M�MݥN��J%��Rxǎ��X�
d���#x�tc^�{C�e't�̴-���$1K�.]:t�!�|��+�j$���b�#��Iv��W��v[����L�K׃,N�*Ձ#�C�ҋ���o�N��������퇿{���\��T<���e�]�7GQ����̓p��	E���w�m:�)�*U{�<��~��j�<19�F=l���Mw�w���`]��{�=7�����Y�Ӿ���h5�<�k_�R����x5�N/rU6�zc���3r�}����a�N;��o�q�:��_��;w����zƂ�$�!-4��[3ױ/P"NUgP�n�_�G7���Ǝ;]Ư�YV"CUbx��Tb�tj�P��|�v��[��6[m_RP�$��o�$=9��B wvvf��������y�qe�P�k�o�眓W'ǟ
��y�8�ط�-OD�_nI�q-ٴ�]�j���{��%	��� rIT���ƜQ 6�iC;y�⥒�yR���a���:���D��lT:b�ӞyvXP��}��)�
P�0��س��<�e��'O�������N@�~۝q����e�eP,�����F�b�IR�iCթ>WP�9KU����w��╫��#Y�z��;����?���>y�$5�y�x5��Ԓǜ�Z�(����1��� ��G��¯�	L��Фs�
bK2�H�`:Vv��w�{�c�S�R66.�+CA�@�=��#�>��6�.�S�1`B�u�]w������׿����X��:
R�1n��ॠ�(=�,��J�q�I�!�D��\tV��3{�ܹs�UG�	6t�z�t��.����E�2n'BVZ*�DRFڭN������;�a���Vz�=��k	�Zk��,��ڎ���X�ցf�z�7L��nۼy���7mݶ��G-�:����~h箛��?��� �Gc�3[5~6Mm��'�a5Li*��)���mв�6}MS���;�U.�$�*��i�T�H�@l*#V� �}��i�MȾ����q���H1�M��������~����&J˫k����;���nw ��N�b�<;)
���^5���a�Jx��z��i5T@"n��-EοN T�֘���i�ONl޺crz��Q����JI(���ġп�3�V��7ttV�ČI�t-�(�&5߬`T�PF��H�4�NM#�
X�mk��J*�h�xQ>�V]T-#S"Q;����v���g���� ��j�䶓g�H�"�t#i��]K��=��]�7dd(t�ڢoV�� 4'�*��d���>T�g'R*��I�й6̭X����Lb�\ZɾgQv���8��뫫�ځ���r�	i�2��p7!N�~�P~��R^����	���>-!-Qd5��gL�~z�B�O�.��EB�3�Z�~&jh&x0�@��P�ڝ9�P P9|���2^��Y�K_�b�R-�\_DeT?L����n����P'����3��b ��T�rCw���k�,g�<�!@�t�]�\M�e���������5�����҂R�'Q0�IW�P��ɥ�P:�_���}ḃIqP�t�m��:6ށ����sqð~����8�殙|��?D��M�o~70�E 3�:A�?��s�a��9������$�,>�dY�#H�8�8Xx"\p˖-��8Y�RY�LY�D�{�)ől�05 �0r��2�8˲�0�X��{x�̱�n��D����T���hMZ-a�K���;��S'�o��)&-�T+4G�X���IWz
������.�]V��e��`�B�5uv���Hu��-�nF��n�q��~��͇?��OB���i8 ��k5�cV*�O����������
j|bt��R�;�T��9�ڞ=�
���̆-;w��`?�Ʒ~�칹������}�d���>��;����9���l�ܦ^�Cw�}���W�z�\��㠍MN$i�X�����E/�O��Gzen����kG_���K��Ae�����uz�2�r�Qڻw/G~��a��ѣ��z�Jq[ j�K�i\�V�/��/BC7�(�|�u�Cu���ġ<`�̄�ǔf��.���f�l�2N����D�~+�p\�
G�ù��~��G2���7l��(���P"�:�����Kk���f��u��2e�.""~���t�ؓ�6�&y����m5��;�uׯ����v��M_~��=�w�s��������ժI��^�2�`�>"���e+����G�0ť/�6����������=y������]�>��Ƕm۴w�����ߛ��0�@�����B�i��*��3TmD�qxx�q`��2�Rix���qlc���'�؃��d!��a�5>�� ��_��`1ul�677wR�'��x�ܳ�>�u��[n���}/63�b���$~��Ru��yt;
�R�ODo�}����裏J3��|�4E�<n��@'b�>F=�[�ɠ@.>��LU�ҍ����Tg���2��������=�Hmd� IfK�O>��Ԇ���Ƒ#g�8}��h�K�����K����Du�޽�ӭfoeuij��u�,����y�����~��=�0�c��������+��Ҟ����A�;���nQ��%W����#'�~T�J������TN���vE�Oc9i##�$3�".�\�'O���q-��D���@_nݠH��ޱ�gwl�z��;�o߼�ޙ_X\__Q�ir�:N.�5;����x-�](�L��IC0@3�EB�Z+�g��^���ڸyk�:���LM?��'��q���33���z���v�p3`��eE+ �;յţ�%V�1b��7�?g�=��,gs�,�kY�~�ȵ~��*�T{�~/�L!�\�@�{�t�&W9$Fd2|��/��� ���K��,2��	�b�+���Qj��������H ��%շedo��~Sx�̮gJ0qTS��V������i�jw`�P/J�* M��'�<��%��k�+ ~L�Hz�n=��������9�7X�[.G*���@��]�4%u�����:4�$�S�u�Rڝ���*�|ܴMu�I���NFYL @H�}x�0D#�"�Ȋ�@!����OҲ�*�Mt�}V��H7�����$K�)��c��k��������
�9�
��hF�
z21Nfi��tc ��!_��MI5�7Y}���yq}������:��y�yޚ�<6k¿lK�;A�t���v ��q}��2���8�={^{�5�l<,~��68�,)��Q{�Y�F�#��11�Irj~!Z���ѮG��A����K�b2�P����$��f��y��8d�4N��h����0#;ي%?M4O-�h�G��A:�c��p��r�L�w�c�$*]�⻁cWC�׿�WG^;
�W��e� i"�~��촨'yM�E1�[�ݹc+>yy�J'����A��#s҈E3[��S�<ǭ?�ɏ'�G�~zq���=U� ��lo۾�Tp}�Ɩ<}���O=U�VU�k� 32{��"������>��}���r�З�go�<{����Uj ��-�ҎM׮[�hήA����W�H2xv#U�)����G���|������������{��)w5�ɕ�ŠUs����vW�k�pe���R:��QSd\-.!��.a�j�0�+�-�{=�$��n�l�v��8�/��"�d�[�`E��G��.R������\"p��ʕ�5�͘�@��,f����-^]x�7��78R��0��ٝ��Z��?�r :�8Z��I�Ht�������c�:D������������mv��~�W�7�mt� ��\��t����/^���3��KJ�}+�BQmڒr7� �M��~j����Uin=��������?��� �Յr�!��8L����7�O�bq!� W�b8��>~�8v5�D����s�I1'�'�~}m��u���B���t�a466R��#��~�i��Q��^w�q8�  ,�3f���8�x��_���*��+k,q5O�S\�X��zÆ 9O=���i�&ƚ��\%#0�M���>��iB�q�R��$��{b�~F�Sns�2�_�M�i�0௛��C�փ ��K/�P(�jr+��R,x~�Fk��ط��C��v���8_^\j5V+e�\F��1u\�=��1l۰]�	�j�B�%�!mÊ����7}E�!���*pH�0�H�
�<R�;}��R��w�Y�0��}(?wă\ϵ�@-ō�f�#6�rB�����0SUB�Ŧ����ƓO>k���vLNO
��Ȯ΋��鎏�LLL�V�W�Z�vw�P�dxʕ�AiVu0۽}GP�W����?������ůÇo��7r�s��:�(�M�DO�����-�F��Z�D����|��O�����4���:�����wO�ҳ� `0X	��"E�EK�JrU��[Nb+?\.�HlW���$�-��Xr�X.I�H�"J�I� �!�`�f�v�����~k��>����������o��}��.��,�E�%È�P�OK�u���N����h�fĆ�N
�#D�����A��u��=�d\\b�t��z/��x� �������α3Ƨ+���!L�$�3w�}q`��&��=����h���~��G��y�
ڒ����kJwD��n�Dj�� �TTR-P.XQ�fh�,�(�W��d�0h	�6%xP�]h�'�W�S�nBJIZ���:B�<�3�+0�I�F1L�f�
: �����)��jK-F��傸7M�%����Pr��@1��b�U����y(��r��I䘍ƌ2�6s�ԅL��F�A�5z��P����?�>Ú��j�e����,Q��X>�Ћ�����O�	ay�"1�O��2���'�%H�@!���p��׬�2�����ѣ-� ��"#���o������b`���3�O�Fm�H����� ���s#����6�ǭi�q�i ӎ�3��/NNN�g�iݬ���HL�!�-@�
̯��c�K;
���K!2>9:*8�5�[vL�}��l.��X2�r1/ɟ�BF�ЁTf�w��x(�^.��+��lF����=v�@�T�h��tPc��L&���gsG��%��ƍ��S��B���f�#�¼d��\�O�r`��2���.^~���?��'.��f�^>y��W��  �B����0�^u����ܷ���ɩ����Ʀx1�@e�^��v�����H��h��8��r��;������.VV�i̙���-�
E)+�9=臃�b�u��w
bw�j�	}�`A^y������}��ǈ@�Ǔ&�@e`!�2k��0�qN�:U(d��G��,`��,�X%�HJ 3����.���e����	�+�JN�9��w�����~����W_}��C8�xf(�-N��ڿ����*�G����,Ѿġ���b�����ݴ?�2ɤ��~d݁B�����w;�����Ҷ0�]ݱ�~�tl��XG�%��%�#�&�f�Sq����*�����C'��x�ƕ��V��_�v���W����(����#�g|lrL8K�t�H�~��� 
=�s颿��7�8���!$�-�E&�'���~�� !0E���`�ٰ^y���V�ˤ���*����`�#n�v��,����1�c1/J�:\���E(j��W^yYZ��r��/�/c
��Դy�[9߀�Μ9��O|����1�/~���o߆p�w���}�Q,"���/��o�֍7�6ba3~�Eȗ��9{�,�]]����+�q R�@��1�C�#�7��CR�#NK���^jm��Ki�q��w���s1����9599>219��`�\��\�ن��~��/�`|b�cO<y����\�i�K�j�|��+�v�U���N9o��fY����0i�$Qﻢ� cC��ːA�z���
K��)։%'.��3��]R��*�\� ��"��&�#EN)�f�s(�]�'�����B�v;R�ۏzipȒ ������'�ޘ��a�ܺ��g�;qOg|t���h�h��L6����:]��Q�R�p��-��}����;8{`?T�8}2��舨�\!Lz��S�W���Y�v��)Cg�`��:qˋ����5���%Nā�#� �?�Iq���5_ٶe6���E��7�C<F��(�`��
�C�e�ňM~dy��0���jC�+�/ً}��$�ӎ�'^��u�r�g��)zA�	C<n�9�RQ\��8x�\&��]C���YB�@��I��#!�V{�SJ��v���A��~�����-��PM j��7�j5��W7������r�A.���Č)�+��Ї܄ب�*����$w��Z�"Q��(�N2�H%�S=���>R�k��'�\�5xA�0�1f^���~ve���R)�����K4�19�f��Jgff�R�X'�߆#�;������I<��L�Ik������i�C|����:/��2n���u�L�&�6T)t6{�����r�0�$'��ԛ�>�A�|�Y��1g�U=LQc�8󼡉�,a�����>Lb�W^yKp�=�@�rV1����1fJ���O� 3 1�@Rl�.��0f(Z 6\w!�f���B|KERaH��(������Gvl:5��퀇�d��E?n<m�DmJ{������7�5�W�^�?h�@>ɹ�k��21y{A��H��r����ہ��/���;[,<rX�8�q�C�{�r��s�����zb�0��_��}�P�l7�#��������FSS3��K_���������K+���Y�M�L�&[��g9^�x��K8�S�W^9�����d�+;�� �	�L���D�
������9y���µB>���}��ُ<�xl�è�jt'�j��^���J>�m����-�$״T*���`�n��+#��^�3{��F��Kv������ke��7ח�ˉ�~|u�f�X��=+�ăl[�n,�sd''�v��>���\�+~��}�͉G�	�%��V��&>)&_�$ڞ6����q��[�����𢡊�&�&�V3���qon!i&�׉%�[2�	N~�FG�O�>-)���w���Vvv���e%��v��\a����p>��j�je�P*��7�C_Lsk�P�&��}X�ё���Z�+���,F�bV+�!�zm���퍥Օ���'�߷�|����[���y�@¥�vC���d�W�G9y�$&��Zz0���]	��M�q-����ֱ�C?�s���y���8����?r�g?���7n���������䨈�B�X�u��L��JA/��� �_|�IF���D���X�$E&�����'�"�C	�~'&s�ݐ�w�Tڈ��1͙'��{�9&�c ��&4��Q�nrT���.�X������?�����V�P�LnI�V��Ti"o�
C�r��={�<���P%@)x(��qT�<8T�8;$��v���1�-&N+"���F�<p�p����F�J�3tL���p#2�1N�lx�<Pm&{�Bo7��0a��s�5���>�b��S����W��t|7�YbPH�F��l����;>����b�f�l��c�(�O r�E���}'���a�{~���/��&U�h
鈐Mba�z����Z�����`����0(ĳ �9>Q�ˮ?�d,�A	�} �\N��<7W)�aR�_�����H\΋Z�%���O� D@���J��zs��O�nl�67z=v7�<W��e��w��&�I��4�B�X$3�
�N?�ruam��X(d�\8�$�V�ך�x�Q�^.�?��ÿ�w~�������h����A��>���$BGVN�~�$�� ��w�	Zۚ���;�lM�d�\���ܩJs��s7J�w��Y�ٗ������\9�$�C�6ԱX�$A(�8fq��~�M2Yi��e�Tr(<.�����/f@",.n�'f��$�O�&=�F�K���:����m0̐��t~�Z�v���߿vv��۷!wf��� ׎�1k�Z��A��Pbj���t��T¥���;��g�5��5��r���_z�I�ʹՔz����D�1Vs�h��L��w�y�*gjj�T�/�����ULE7E94. 7�`�0�o��������Ȏ��u����� �3�"��a7r�\��a3-�M�~�a<au3o��qk(H�N ���NbFr`�S9�&���c�ٕ�<;$ ���u݄��z�]w�����1���W�wd�Y�6��K�$Ǜ��1�$ "17��u�}�] �a6Ȧ�;���e�'��?cH�9ؓgΜy��i3Gd���*�%�!:b7@\�i��\� >�`�ͩdzZ٨Umb���.����X���H.�����5��ڱ��$�"s�0��d�u��n۳�е�������g'J�P����?������7/^̾��jhM�L�������q�7n�Wj=� ,�R��m<v�W̃�´`-��>C��htz]=���@�ׯ�ӟ�Wʽ 6V`GA�Ve�J�X|��1�O|�f��j�� 3ha���/�[�q�̽��y)c5��:26�z,�3,�����ɾ�z��4��䖒������e*6w�M���c�#��ŋ��xh��gV�l k���h4��[,c�J�{��˹w�����j8cb2%:GW�!��0�����a�`&1�'?�q��LN\38���Z}6��h^\\��c�� PD0�>$�Mɀvd��h�#㦘���e��)_�t����Ȱ��A/ի��
������ؠ<O����f�%m��+����ɭ��Z��Wx��.���8�r�|F#)Ȅ�/��pme�T�h�H�I�`*G�'��օ,����k�N�>��k�����|�\���GE��q��G`^�����W���sM��+�Ȇ�����np���_�җ~���\_[�r�l�t��qh�y�$�R�������� ������3g��v�ay[9��'�Ǥr�^��zAM�Q�N��L��Q���J7k�D��,��94QYqi��
v/tG�Zh)?�u`	�,d�f�����BbΗ<��v?�F�~{sk�\.9R�a�?%#�$��v.�k����'#�������(J��+�5q�K�fk����O}�����=��'���0��m<P�V&�&[R�'ͦ;����o|���+7n^��j�~�X�泹|F#i�<y�.	���Zh�Æ%��~�[AXȗ�&���Z���l�8M���g�6�,�������8��˖7�۽���=������'������Q�OH�m�rKe����Tȉq��r�3D��W��:��%Y��o��ִųS��]o�Oދ�]hb��϶�"iH�VEbla�"w]b!�|�+�zm'p#���ʶ��7�;�V�8Q��b7��>;����t/��h��Ug�*����D&cr�0Wι^ގur[&�O�H���
2�e�U �8��ǵ����Bc~~2���l'ꬭ�t6��J9ͦ�^��ӕB��g�.D/�j�N�Ŭ�(���vU�S+�2^�
@Y�ӎ1|I;a(`�..��0��f8�Zfj2,9 Ff���F��9T�I�~�L�Rǔ��U���+o���o�A!>�_��25XldD`Cr- ����������7r=�Y0r���8�@�OǛ� l�M��3��*{��3��ܿ�bF���W�+�������q��� HxX|��s�������ø�ٳg�܊a�pq ordK+�e�"|��B)C�β����U�?�-�	5�h��Ծ+i�����LJ�aT��*4}���Y	�]D�F�0>`;65\�h6��bzY/C�tB��3��R6�u�Lvemub���A��}��쁹}ۛ����C77�pV0�7o/�/�>y����������jw�ff|�b?ǰx ��c�a��x�;X&H���e��03��j�x��;���������r�B'P$jw�d�4��7۝�����/~��R%$-�ğ�۲�������~�_�oJ/�90�´)6t/��'�x���\.�����wO�;J6��1��BS��5�z��,�.}+�b�����ٜe���|����1b�m���cbT���+HMi�z���9T���:�?1/HTa���3��.B���h��?��C,�j{��c���6��,�Lh��rzz����ggf��xCL���Yl1%�9r��eb�\���+AHՌ�%o� ��_�yq�8��{�c;j��|^�h�Yq5H��^z�^��w߽��g3��i�I�;8�����G����(F,i=�Ȝ�[���d@�������^w�T�0x��Q��f��
sf�����1��C���)�U(�{�U��lIG�w1�d��?�|���w�A�{R5�*J��u0s�}<����=���7N����ԡ�!�{U���M���:C7����IQ���cF��uw���I��w��_X�&b��(�!y` �R)����߹���AY�l�$����pŢ�2���D ����1Z��i��(�GLU�u���B�z�Ȅ؞l�8(�O~������<f;/s1�Ӧ)	�Y��	�?9�+�: ����#{������?��(������fB;��ʥ�����j�����^�y�e��"�CI��@n6'�P�f�\��:���:B:,�~y;�:��[�R4���[Y؆x�v������ձ��������c���e?�kKX��1Ϗ�Y;�!�؃ړ�@FH���u���h]��f��~�e�z���P�'��рM�9"��A�'}�'c{V�O���=�}w��T/?k��9��(dWPFM���hn��jւ�fy/�B+H���s�=�*����O2�g��
$�F/��i̙!/F>�Yd������>BI�g#N��:I�"��������i L-��N�#�`���<��8�Q�P�1�B���Q���{�yʵf�s�4Oy�bg!�h��Ԡ�X��| 6�����I@tA��00�$,���G��b�LW#;�Aȁi�5l`��Yc x���i��id#���j^���JS˩0�v��f0���x^��ih�G�Y��)|�z5X9x@6�)�_�3��^�~p����q�X�y6�Ό\�g�!�3��]BA<[bH 73����믿΅#�*����*�u��dY��U41_N���#�J:M�A��߹th�!8��
$sA��Pf��`W�_iȹ��|���j9=p�޹}�a��jom�[�c�Z�`H����Z[����fml�P*?yW�X~��Ͻ���<����tG=87=;��o]���;s�ޑ��j���)��L�0�7��)���"�ֶ�[�ǎ{��O_��Wο&u&������(!�[Q����p{~~�vk����O��/~1�Ϳ���޾��ONJ�/�+<�裿��������ko�~����#5Q�m�V���x�{쉷.]��×,��^�IzP��bx�$8#�*]|���%�ޜG."�֨Z͓Y�=��ƛ�j���8�nQ""̑4~_M��V�3k����`݁��*��n�}��R�0��^��w� N+NS����!��q~����&��#��!w#+��tǢ$i[f X�=�ó�Ybx����lf4��%z +�W�1v���{_���ę"~��U�BD��?��
ͳ�d���nͭN� 9Kƿ NI�d��b�A��\�2ݖBÐ^3I����"6� �K�\�t�����,����]���W��2����}P�(���Q ��$��e$�2Z՗~#{��
3���cd���������	�6,��k����JH��Hu����X�n3MbTt�$P?�yn�1T�k-q��vԠ���R��_!U��H-�~�ra�Bg���k�K%�i���r{a�X����e�	�_�����-kqE�n�P��%toe\��t����I��S�yߺm�3̳��IH[v����_�;���'�~��Tla�J:�V}��gbRFF���^?@��z-(қ7�7ַ`!W�޾}��Z����{n�Ri�/�Z�������8����d���@VM5}���
�$S̎��t��V�-}�4t�6��oI6���PZ�;�N����=S���w<;ʹ;����r}|�SIx~��0��;�U;����L,�]���i���섀pLa�V��K�l{�yՀO�$V��o-�ԁ�c����D%��^�-V5�.ն�1��N>�،`7°�|e�z-3R+G���0A��v���7o�;1Rb4YTc�ım���e>ÈT#�F�O�f�1�L׎�el �j�#����L��Z}�5��̗�z����:z�ƭ+�_�����>�F��v���a<G%����X�YA�fhN��7xw
J�`�f������!���Y
�l�XEs�Ӿ:�� ���Z����p������	+Q�h���8$-�Tq�	�7�
wثp���hW�ͳ'KV���X���@ꌆ�!X����P��`���l��M��|X�J��b��b���bq0�/�D
f�,�%��NdE5��e�,}����=�}�����	e�a�U9{+w���=��*�5�����6�*3J���d�!Dݨ��ɵ���y�����1e����h�4�+����0��0�?��Z9d.Aq���̗�N�c��^{yiy>����:|4���Z�ur��V;<p�%e��́��m���p�쁹C�3�W/_��2��Q&y��`�w޹\��f�*��Ҧ�Z�,����מ={8���^�3��\���=zxnvv����/�B��^����?{�=��C�LO���kk�~/[(f{�g>�b�r�����?���˫��f���­�\��?��|���8�ͯ]Z�\�B��ŷ޹zy��d�>�3����>渹�齳��j���d,�T�0=��V��*��A��w�L;��U4q��\S�Sz�A�.D�x6h��Ҁ��;S���T�(!} ���$Cd$�FAi�T>)�4� �U��*>|�5-i���[����6�N����(޿uK:D�ݻ�(���8��Y��w��Sy��������6p��b��p�S3����#LA�Ӿ��^,�� YY[��l���C���Kwv�0Q.U���Up���2=�,��v����^��z9O*��!IZ��t��_1�VN���l�tqqq�7���WV�QIh�$��o�.Q7����,���N��&��:�9,#�0ȷ=�{>�я6��vI�2���t~Q��;DS��𘔪�FAu�)��UOǝtg��JM�����~����f�h�v�zK)lw��)�R�>�6Є�/ޚ��K�z
&�Y(H8���΋�6�n?�� �jؖ%7��JZGv~��ۆi�\�D�ؒ��~'�[.�l�a:K^�cb��|��z`���ri�c'�R�cO��K_����Ƿ~��Mn=�����?��Z�h�3��З!��V�Mo޸}��Ml�����k�:�Tmo7�?D�+t{��K�AH��>��Ry�.�RQZ2lw��[���'���D����Ɔ�Fà_.���@��~�㏏U�f��
�|��-{)0�*�M���� �#��>��Di^�jz�d�T}|���H<����p;ͳ�O)�yJg)�3\��E�ƍ��4���,-D��Q��0	�=��`�/��'6���$
���'�:��=sq��m�c�ƀ v�9v���y��lW�'�\M�6�W!�q���776�`��4{�ٜ'��%�6?�?��ԫ��A*�)uȸ��[�����.iXB��>����Ri�"�pM�*��\MuS�Ӡ4y��b�J��*��aS����xG� %뤍����7�n}"\Y���a3��^7~,�	9-�d`��3��鎖=�
ۼ�;�\}X~^�X�*�%(�Lg3�S�X�Ġg��	l̑#Q�.�I�dl�E�c�:�HB@�Ó�����S�jQ1퐭��6�.LV���&�XL����$�Qz����USg:뉓�.O�h� ��
(	�v����d�8Q(�*5��	���A�z{��%4}��ͭL>�/��|��W^9�G���O�:�Pl���ʥ쾑�)7�o�ڣŊ��YQ�͗���^��R��nUGF�$^YYe�+@�R�G�-�C��GnC{aa��hI��G ��W���K����o���?�䷾�ggϞ�|����s�*X�O<�؃���0b��H_�r�(��Wη[���k7�o\�=19+@hzf�6:���o��|���u+�y聇~$�/}���.�^�;'�ԹȽDf܂mF8~�K�Ƣ�G�Cw8S.�����ZɰT��p��T��\,�����w%��%gv�N�4�LMMa�3z*�>�+9N���ˬ\�c��Gu��Ci�Z�ZU����J���Ȅ�����NUI�<dF1 ��ѽv�w��Ë���idv���I�I��t�����2/t�޹r�v���Y�D�Z�X�BSd���;ݒ�_�~���"LL@?�ƹr�b��B{�x%�?f�X3VA��eG''�ՙ�G�Ϟ<��܏��<�ؓ���͛�p�PS��4��.��?��I�@����~����k���?��Oc�蠃�V�s����Wq)EӅ0@)2��cMRC��^+r�M\��']o�0;?W�)D�*�g���?=o�[S����S:y/��YnDeͧ���t偀�L>W�_DL�[����W(�ayml4�����DAxKjX���~���cBVn��f;��Y	BZ���2�~�,_�uL���_�D�z�����ʯ��c'Ӫ�)\��_��_��>�=�m�T�8��W_YY1�$�{f�9r��7ۭ.����v�ۧ��z$`�t��Èy��+�A�n����{��#O���_�x�����gN��n�v�\~�ٸv��$���&c�v���z�ɺ��ՍkW�:v����r�x��Z[����g}�y~k�m���qf�c�������{>����@�f�-׎��P��L�wʅR1�}@���F�e%�Y�U��H.Ke)Է�J��nP%�<�	�D�P8���8r��Y_��;�,4gi�<>36R��7�W� g.F^���+�/��M<N�Ս�FI?"�� �K�v������d��2�����Sʗ�3�1��/^�tI�����/.��K�!�#�4�)�i�3C�֒erP���0��2��3/�=�[��ڞ���D��]��
��Z��ԕ�WS�5��$+�	�qT��(MƐ�vB��V�0<"N�R��F�!�^j��й�a�'%��kV�Ћ��Ж��m��N�&�F'.R�ĩ�!b143mh�r8�����9xTfJ���u��o�v�fe�l{��R�j�Mi�Ig
I���rU��i��W[Aa����S8���jr&���qL!�4ǹ���eNx�H��O��8�ǔX��X�7Ω���o��L�O���}��x��t�5��V�z���ɜ��Gǧqd� r�́�C�/��9Υ'{̊�nO�����=3�ݱc��p������)_�ۦ�Ǵح-�af,�|qq	r�^/oo5�ݿ����}��յ�5�?X�ׯ/���g�}�3���_��1:>.ʒ H�q�ԩ�Wo�۷ou�s,�С#������G��VW�n�^�b��g�T��VZ���v�ZZ_]����v��/�cB譡�݁�b�!�cI�򠯝���%
�X8�k�~�3>1J��y�lQ��,����1@�VZ9�ݴ�Gm\5|@H������u������+��"�3��-���I�ٱջ���@Hy�I��R+c.�:׉�_aiLZ��O�%ó���!���@�,��N٢����D�w٦Fc��w_FԱ��zU�R�%�'��n�^��~�=:M�(��;��lmB���3�mzY�<���t���;y�����It�T39�I�/N���®6�ݵt���7Md ��r꟢pNW�07[�Ꝁو�����l���_����ӧ��? ��[��������]xffS��CA��߆����?�ԧ>�J!�|.,,h�����nE��T��;ibM�ФS]w�����	ce����pVC��{ҙp0�vܹ��n7[/�{mv���'��5�@{f��f�x��R��^��7.s�h��e�� (�+��k���^�����'']��v��rl�!%5ζ+IG`�޽&N��a� +��Lҍ��J�[�XǏ���>{�=���/����?��7����W�^:;>6��l�{��fr�nF}C��kcc#&{"6��J�B�տ���FqH�X#��ɑ-����R�v��rA���2��>ί���{����q��Q���s+��0�N�T\�Vkcؘ;^�V+z��卭��ŷߺ�`�Խ��՝4�!�1ű=��/����!��` d�'�'��=���[�W~��O�����No��꭮mM����dy9��xF�K#�t��&�����f����� }�2L�)�z��&bw��F����/��Y�"�@��x�m��-�<;%u �p���zs���ڳ��J��Ey���0
��L�\,K���$��_9,Dӹm� �����043Υ����.N�# �gz
{�E���	�sޠ����������w7NLH�N϶���s�Lm��괉L�4\%�V�,�m�� ���D ���)d�S�S?���X�A��$.9�w�����Ҭ�(h7�R�}2^A0�MB�Y�Z1B�_z�(��)�Q��i1�lT�ʃ7��	�����$�"za!�"L"�F�I�FN$�}ʮCM�E��6�ق��j�6���!V���3��p�</��.�V[�*B`#&(l��+<�48ܚ���hz���̈́�9� �{YD��ؚvVamA�n<.A�����tj����҆��$d���%���9�ܕ|akkK�"�$�@bS�>�t�T������t���~��_����_�η����l�<Z�<r'��5�nu
�2�����r%N������~gscc�����]�z���f������vcuy��8�Q��)��-d�wz~������v/��3=5&o#��wXN�ŋ׺��t��Ѻ��[�W�\�*�������ڦ�sZ��v�U(���v�1R(���`�<���^�����=J:aw{s�fsK�y�5������L#/L2l��l&��5�m�GyA�^ �Bf�UP�)I��v�	�����^�\PcZ� ��4"2�Iu�����k7����WH��+��2������	�ˈl-�1�t1���J����<P��\��#a=�宻�J�̓2�*�+_6��g�㰪���(�Y�D���1����J��.g�D�*�a�����I��{R�� v����L3��R^z������O���-߾%��R�a�t,{�v�b�b٢�aP�����ƠB(�dl+���$Lb�I�t��X�N�X��N&�}����m&hF�h3]E�v��,�h�<SS��v�EYAwd�2j�������o�߸p��������#��~���_��_������RP�ح[�^~��g���d����ƙ.�|T�Ud�a:�#Ŭǔ�.})�Ji�0)w�xA�o���i�N�� ��^��_y�܅L6�wړ�c�>���?��ğ�$�)߸q�ܹW^9w�ܹ���i4;�$����5ǎ~���c�J�z�'k��
n 7^x{�v�2rum!�v��l�9�w����c�>���*��.������o��o�ƹ����^W8��Ğ��#;�|��e�h<�ɓ'!���V�9uK	����}��|E�?4@'?p�bӜ�1�1;����y��._~��s/8���������x�V�b'����^f~i����w;��,��1��n��,o.�n7���������x���} �RE}�'K�A]���D�ۘ:<��_��_������ŷ��_ZY�v{���{9����[P���1��B�߱� E���6S�T5�)�^̒��}���QlG��`hsȡ)�1!E�FaF:�[���NI�E����Kؚ��[�v/�/JU����R6��I��/
�{��m���7��7]��+����V�!,@=�|7���-�j��|;KQ&���R9�J�B�o9��SLHѵMA^b�m+��`�ž�xB�O��G�o%�d�V���S���|�<��[6�v߳2%�N\�'�*)�HX9�;�c5;LC���v��bN;ݞ��뎌�M�MOL��� ���V#)䋥:}��$JZ��E4(��^d��q�Ǵ��I��i�R�7
��]N\A�CiK��++7�W�Rv���#Mp��	e7�DJ�A��&��ZO����6�\��h��r���$l'��9l%+W,DhA�=�y;-�UxF��I�4+�)p�~����+�9�ɠ����|h��j��!]D���_�0��q~��f�>�X�L�!MAf-n��T�u�U��0F�Qq�	W8�Z���*���L�+��ނWK�'�X�~�j
����dI�
��%���_�W77Z�����n��}��~uz�Y��~/#N����d��v�7�9y�O}
�����ypz|bk����.i|leeifzo������.��#{���ة{Na�8�K�o޸����+c����� ���#�Kbd��ZZ������>�q��,���39��kK����Dw�k#���v���շ�z�2Z���|�|������a��i)�'?����ϟ{���>��I�I��h���+�SI���c�\fb�Z-HgA�4�҇4:�yx���=�j�yyI�r2��� �Jذ��~��q�j��;5r�����\�����ˋ�bJl����WLc��qa�Z������ǎ�8z�me�a��[�o���k@���� ����*V��ʣLr��v������[K�Zn����&�"��\��LX�[�j�N(X���M�2~���׳���ͻ0E���J���v��5Z���w��}���g����1�77����;ҜN<�a�V��\�jo����+�]ycec}td���Z�ٶ-:(w�<�:d ��6�qj�*��RΛ�<������DV��������p���z�w�yGx�#�})Vt,C��X'N�u��q�M�bh[B	�$o�����\�d;amnl�o,��/A݈�,�!$�HMZ4,��$T�7Z�*I4�P����e��l7o^g�k��a7\^�\Z�8t�D��H`Hy�/^�|�[���s�=�\>\gӼ�|H�Gٞ={��?�G�����}�ʕ+�<�̑#G�������bmg��r&����Ԗ�*6��_�vD����W�S���S�=��a���')�W�NF�ɮ��V׃E	\�%�s3#$����?���a̐e�/���/��Q�|�ES�i:�1�����y����l�T2i��t�Z �,��3�����j��]���r�>����S 6�'�rV&���L1s���\~�P�{����W��+_y�싕b1��R~m�k��H�<��:n ���C�o�߀yyp�o\[��h m4�Y4�9���;��y��	�&�c��t�H����܍���[oByU�#���7;����2�����v�!�jou�~'qi�����z��c}�$3c���i�N�����!�Er%Ҧw 229I:?q�����8k�$s��G�kkKQ���Ǯ���'n�Bp�]H��:����؆�U(M��H2��C'��L.�˴�BF(��ו�s��~��-�:�K��lz�S*g}�W�"aז���N�Y)�m���]�0��f��p�C(�n�}I������Z��5�F��U��$��,�l���]+����D�=��*�m�\5z?w%�p$T�;�^[���$���[ �`�9&
��Iy��Ќ��]�2�Ww��Hj8R���r��Q���J��h�\�>i�ku��1�:�iM�G����Ě�:b3�j"3�C!�IShD[Yy��M!�9~�v�����L��hʓ\N�ԝ�..���^Jv��?i�R�+�8��� ܚp��vZD�`�B]5�h)|���}�.B�P��څDM|.��j��..ux���0��KA�])�:NN�f�i��B���J����ឦ�W?\�6��LZ7��� Y���@�aX����8���&��)o�uI����Xz1��f{yy�����ɍ��f����'GjՕ��7n�Ll/Jb�*�d"������)ȳ~ܼ1������[~�42R�����+�۰2~�a���{�=��S_�������ZY�ƨ8��5��9s���=�|n���[��Z�͛��?p���!
&&�WW6�Ϳ�ͳg_����6��8��ϟ�_�
�(��\��])?{����;r�d�P�F�"St���g�9��"����T%.��ԔI�2��~��k��7��K��L��Y]]���d�p�f��A�i�kR,���̕bռ��p]��h���^}����]�a#��?���y_/2�'d���q}�����v���Lp���|ĺ9I#����2��R�`��	���fI<H�3������H����N
DibS�ο�@�P����$f����i>p�G�������tw�2��mp���S�N���:f��,޿z�������9���a�)�^5<F��r��+b���ߙvK�����x�ɱ7���&j�HO�i}�V�g#�W7�P}Pb�~��9��?��?b�P�̉�	�.�={�����<6��|�kt`�:�!�����5{ ,�v�>�(����gM&��WS���I8*v�f�%uu�>;���;�<ӽ�i��n��a�.:�v���i�p�S�������g?�ٟ�ٟ��������n�j"剉XV�~9���-�� 1��f��{��쬓ĝv7�5+_,����/�H��Ӡ�8�{�I�����Yn�*�9�3d�Ϲ������p�u��F��%���BI�a1m�?:2	,���5i���$����+�s��۩(dq0���^��+����'O/�rt�r�@:Z���ݤ�lݞ��}�6f�����މ��C��\ZZ����)�/�GK�"�9��,���_��6������+	���z�����n��,��ܖ�.����`U���\1����a+��cG�:^6�#c]��C��s�T�׫B}�m��m�(XNEׁ���8�j�����L6b�~��fsy�����p�'F'z]���T�$[��RQ����h�^��8�G^&��\!��Pn*4��QN�!]��C 4L.��e>6E�@�5	�Z�r�9��a�;��� ��nM��gh\k`��M����@�Mϖ�N��ZZߦ�a %��R0�5ZJ��}�hA�2Hכj�R~�}�t��7�4K�����0z���HǠ"X+vh�kX_kޚ��NP�ړb[�ﴵS��tT9,MI���oY�~y4x/�b��lZ�Zk����*m�Ri��t�7q���j %��R챫"��4{�;'�e����K��r`�#�P0��2���
ZT#�9�8~�X4�uJ����cZ���ȐOyc9K�
H� ^+����0/M��H�?�w�^�kv]/�S�x8��n����ѱ��ٝʕa-��m�߾�ˋm.E��B�Ӷ%�o�-�b�077��W�W�^k4�s��w��~���1�:�er��[ׯ��g��ݻ�T��
rN�����[^^��޻��?��O~��o_|�/����׶۝^7XY]�;;�˿�7{���ş�NL�E��?���͊���C��$�x��-����܅1À�{���ν���7K�zl9����Ravv�K�+d�l�w�XU�u��*/��/C	gs�*��SSG���c�^�4�]�U1(m[̢0��ZZZ�������w@�e��5���#��0N��dr�?� :���$��m9�)'N�̛M[BC���ZA��0]h,F����f�T�98�vCz�%�a���� �Xj�6��*�hD��L�+:� ��Ż��x��1��ϸ�q"�;�...rf`�abi �n޼�o�Ml�W_}ψ�4�!��A��G�N@�p�Eq@A*�VFF���AE^�z��_Y�4E�ۮ�:iє�?�+YB�U��������И0��|m�p�����;���*p��+�����d`�t����6PC�L\�-������I�K���*� dk/lQ��;F&ڥ �^�}�>)i���3]C��(m ��`�2>�=��o~��G>�kPG��ǍLLRcSa�k����k����ϑ�/�j#ͶЁ:^ƕ�Soee����~�pHg\�Jޓ}~g3씖%�\�SW��0�Y���QY�N�6��Rq||l}k��^ƣ�rR�WF��d����0�����7�5� &aX�-�����v-_�p��Ņ��7�Y����ajL�a�Fb�A�v����ޜ����=|h_�632V/�w��^��ٳ�C��c�Ю|�t9���m��=��Z��EN�j�s�L����ne�Zg\�/Ȁ�<gfj�^��q�P��Gk�}i�ṀCIƎ�� l~�<ڶ�q���P�K�PvI蹙b��9�n�!��8��W�Dtf�a$76��ڝ�_(zV�qm�W�P�E�e��I䄏}9YH�Rz�Y��D����lw[�9ϪԼFݏ�9)9�wc_H?�2c!�w�;
���+E���Z�$��nV�g�*nH*}��v�D�Hl�;AӢ�s�ѱ�$�loo��FfҮ2�~���v����jM��l�WIU�@�D�iˮ�4L9x�U��`�¦��H��v1��%����CM��I�b^5h:�ߢh���$.���k��^��(w3o��j�s��r��T�h'%:�J�i�:F��5rE��qe�U��ڶ���A(�L6�s���}s�Z�D;��*zg�@���4��a:�H
�T���P5��;q�q�ڷW���RBXݴ4����ǎc)N���c��.RnZ��䘕�Vsl����me��L�Ă�0�U*�m�^^q�����$J��ð�"�2F<FK���m4�MVd�Z��u�]n�=��ٷ޾T���������rI�Ǿ��o\�x��jLG�崹�����#c�q��X!��ڳo�G�������'���/�|��ܸq#r�u?�T{�������e�=ӏ~�L L "��#�X�R]\��B����~�c������&;6�Vq�k�;|a���<KƩ��rIȯ���ra֔��r�3:>1֐����-p�n�:���?�!����U��+��ap���J��!��Y�0x�8�L]M>�6��<kX,���꛱�	�#��}Z��p���Ҹ~�G�++Pi�>֣�;55����Z��I��	Y|v��%��u +���7[l�u��f3���] l�֨j��J��)�@���� �#�<��r��Y�I��p���.I~���~���->��Nej9�>�$�����+O�LE�v�^?M���łҬkj�R����h��ǣ�`�/\��m���{���YMĢP����u�1ª��G�4�1�k5��-�jeʹ3<�$�g�*��q�Y�%��c�o��.Ji��R�w��k�
��ew'C	Nf������$x��G}�ԩS&��'$ñ'�̀��0�p#�|��w��.]�{��}�oU���o5��l&;ط���r�;P��������u,_(�r���#S�	q��O^��֫�^���KU�(�C{��0��csQ�-..mnlC�3�������!�#/q "���n-�V+����#�%&����LWN>�����#��tm��Y8�^.k��ll[�� ��;������$�z F@��n}b�C���@H�4C����Z�چq#٩�~3L��>�V�w���m����T�gE},Syt�:R�d�N��zv�X���� ���H�`��c+� p#ȑ�'�	���c{Ya��`Y�8L�%> .���4�xF�\���jDQfd��	�#�"��g�(�>�J;a��C��<��R��Tjeǎ��A�	����W��f���#�ω?JN���V~w��I��X)v�oB�V h7H3�&B+y_��4U�e��a�N�ѹ�����r�>d�Ԃ����K;���"P�B٤��i�Eň6S���-��6����敕U��hht*2S����B��F*p�oY��7���$x�2�8N���@��)ԊR>=���=��%7K�t��Nu�ҭ'�.���!l�ސ�Sry����s��cʘ��Dz�4d� P�=h�ҦIO�.�I��D���Y���ʁ�SL�=V�+i{:�Q���P�f ���g'�.�33i�Ddn�ڿy�&tmG�ƶ�%�E/��QO�I�Z���Ķ[�]]Y*�=?��U�,���F�D�	�巻^��ؒ�
ʅ����0�~�>*�#��V�e��^�r�ܹWx9��E�Gmll(�1�_�п�;�c%�����핣G�����Hdy�R��ʛu�z��e����ݿ��SO�������������k�n|�����/~�K_�t�������J���U���ko���3���x쑾���mlkǞ�T�d��tdX"���H��%�D�WV����7�..��)y�Pu(HYw!�$�2#i>1E�i��]#Z��5Bϡ��2��.W��ȷL�VYXX�e�`�Pɔ�t�u1�l%�\a��l�cǎI#�^��5���piI�Y'�eԢ�{�,X__�}��a`Xޅ|�k�=h([aHS�Mɑ���?1L���<y����;�.]�ysޜD��C�a���X#|(�̙3�_{�F�EI�4��W����0��8��(B��~�R����c6���j���| ��_:U)T�I� ����׉3�\{��R��lH�$X�X�}��MNN�3��Ќ�@K+�y(P�k2�cް���U&!&���I�yz5�8�N�����0.�V+����jW�6h�b;�T��XN;�v:"��f���hr���[ �L�e�c�d�B!W(�\�#+�35�������������K�"���r�x%ʱ���=�ߚ-f�n�����sa �|�,��NݍɊl/��j5��SO���޼�p�ːP�܁t���cGO@daoܸ�������Z9��R�^Q"F�-H�f�56>9>9���O��i�T�Ąl63�z[����0�� � P�w7w�g'�1�!1�W��&���1�Il$���bc`d�\��Ŗ���|� ��Ql��xq� ��n`!�4���BK+1I`��� �����v�D"#�F��+��9;6�e�T,��ڽ�4��W`(v;����r�H�긹N;hwa�8��z��i�z}��z�l!r�!Y�i ����В��V��q�0�&q7�ڮ��ٽ�&��_oZ�-)Y
}��r�~��NS~uޛ0�LAÞ�x���>o��	С{þ�R�G�e'�zR )���\I��N;�)���Z�R�����(ҥ,�\��|��BU�T�|�7��M&�����e�;�k��ItZdO�I�@�:�ԗ��;���<�s����Ly�ԕ�Nd���q��x�V#E||%���|:od��VH�NN=�j�p���TMCZ�6�x�e�S�Ѽ���ZG��(ϵb'�Pk�ŮT�װ��T�.��`�����]�$�LTs��ɵ�VA�F��BJϕbfx�"�$�٨%v�8k�i���d�*'���u�o��+�c`���ϭ7Za$��W�6������߇���2�n�]1U� [p39���C����t�1�d���7_*�{TF��l���#/NF�c�6����7�+��z��g��B�R�e�����T�R�/����,L
�����/��_��'��e_}��f������������o����_��ɉ�'O�8q��+�N��"��ԖÒ;r�XgϞ��69�9ֻ2$uu��p$r�</�@�\(5xM��*x9+� ƛ���ƺ9}Ł!e���u�O�4	!1�dT��ilњ�`4:ѡ~x��.�zyy�a"BZ1�.��V2�}��Ց�bI�־�}�v{�Q�kh���?��w��b�J�eT{���/^|s~�����7�����?�'� k�q=���YW�t��򞛛3���"�zR3���R��h`�ac�{�x��^z���,�g�&��)��,��W_}�w4u���i�0��N�U�M������g>/tMn�_J����cgM�ޟ8"�t�I�Sv���;C�`<.\`Y��U�<��,�}�c��9z�(��1�G	���0��K	��a��6���i{V2��>;��a?�H`Y�
[]�x�M�Y����wU��T�t�]�M��Ki�qW]�G��Ȣ�	� B����$�s4=�iO�2LǍ��e�ʒ]�u߾n����vK岗	�7�x�M�r9I���8'8��S�zg�6���(	�Ԋ�G}��3�c�\��V�T�Z0�0�i_<`��̖�����w��6VV�VWW!��ɂ\3�	R1	�`�����T�1�8	�n�mn�����{ؐ�ӗ2q�Բi0岐V�,��i�����<ł�A�G��!�Nql
�aJzV,	�|�Tɋ��� <���Jmr�499Q���}��N;t����&L|��V�P'�eY���꛸����:⫰�@H��$�A7����9���s�+-��.�IK��b;
���$�b&W�zŜ��i��������K� �v!_�#���Q/ ��Ts�"�O�������Doe_|n���NR��;N`TQ��0�F����qL�<8TH.�`�um�г�Zm'�2.󎼞o��vq%���:D;IP��M��+E��[[�<���֔��K����DmM[��#ݷZ��~D�E��z_�3$QP2e9��X��j��`�X=�dV:�`�bb�E�:�ҹ��RZN�����x���}S10ύj@��tf��3)=vć��HY�p�}ͣ#t��]�[�)di�A���]D�Ѥ�D�1u�jtKے*�ђ!��Lt:�ꆶ)������)N/�f�BA�8�}0t��i���������Ҝ����p
k�-}|�����&��0]{OGĎ_a��Ki���泹$���ZJi�����֦�6�NR�W�@�۷����a�ۇ�,VF���ϕ�l�kK6�#e����\	#���Z\^�u�&&Q���US�d�H�#�ET�f�kHC�С9)�.���0���L��,��qBa�	��X�8�x����������~�k69���Z�W*#�'���?����_����Z�I�_/��Ղ�XYZ���q��0�9<Ԙ6;ٶRMNT+AX��ɉ����~෻�l��x�`����WH_v�)a��~8|�����.��]/���!1��ӟ�LqwL,5ʄ@����;��kJ��3g�@��;�.�<� ��ٕ�X��~.9�Rh
,�k���|�byy���_��6��H\(]a�s��م2�a0c�>��Ǐ-��zm;�"T�C��]��i�H��i<�4���޽{a�c��;wv����p�p��q�ӧOc�ϟ?D�9U7-ţv$7s�ӗ�,��)��C0,;�y�����k�zWN�.���BD�m�@	�m� �i���i0�ex1"���I��.�����jw��
s���U ���^�#q L�` �JMeo:R�>5�;�L��O����Y����M�tA`�΁���j�ܭa`M���|��8=AdX�x��6L�]!�cw2z�]XQ�HPr��q�׼����a�8ؙRM�w�b��C�>���ֿ�M.,4�|�V�<�~����̖�`�B�"$�3s��d\`0��.�G^661�k���I�
�B��n6�(6,��q��P4 B�Bn���vqw�����fC�w Vr�#B����BΎ29��b!�w���7�L/�u��B��効>]��;upnf��D�+�����N9��{쳜�p����fGj�r��B	sF�3I�F�(VFh3aHX�j��V'���)LV��W�2�&14J͂0ȱ�) �u�Պd~g�~���t��������*0��ʔ����.-̿��������J7�"ۉ� �+���@��sv6�T�X�u�趁��n ��-I�jl�~�)���QQ(��.�.��t���F�%���irݮlZ����z�-��YiK5���D�j�LLL�����*-M�b����$�b�R�Z���Z����֠G�)��hB�&���[�j(�=yئ��lT�����9L� N���e��>8#9ip��fC")']��[���N���	Q�\:�(���b_dZؓfn�$r���S��d<8�3g��"�t�Y�J5�5�e�Ф5U�W<
�4��oik&ڗZ��5!�1>ŝ��	���#Lh�����A�|n��s��um�S�F�j��=�����ȩ����A؛����oZ�67���,Ȯ���_�s"���<� 'p&M��,ږ[vے����P������迮����h�>�QQ���].�˚eQ"E�#�y@"�L�<��ν�Y�\$ U�O��R��w�瞳�^{X{94%q|����0���N�^+���Zmuez_MNNb���W�-�t�(��5=:!7^�n�2�k��6<4�p�>�X["�=�Z�����S��V��\^^ś�ᭇپkw�������f3yH@��;s��,m5�\�^rg��u�N�jfb�ԑ��[�$��I&��y�)/a�����w_q
�۾��Ȑ����~Y�y"��<���f�.s �RO���D�h���F:4�`�3���]<��Hþ8t�Ю]�0��J�T.'b���f�;ᮇ���+/-`�*���]XҩH�ХE+EP�]]=��
�d��ٹ�m�LV<���홛��{w���M�HrS�a*���r��U�7�x}��] !8�����ၸ
�SŤ��tF�ޭt��d��^׮]$f7d��У��i��<��=u�ԕ+W�V��8�����D�8�0"�����f�(�uܰ��8�æ
���fO��_:����>��5�|� �Xu�ᰣ����������}��	:�tC�t9�Q�b�������ې�hA��J�p4��v������Kg��)JG2Ӳ4�I���CJsWh�#��fo/��h����j�F��G&��3�gO��Mǲ��Sݠ--yb9�J��!�a���Vv�q��33��|��&�����?=�_,�3Y �t�,-b> ]��u�o�>44D_�Եk�K��t&��^�e-o�Z�I�ƛ�O�W�R�*����	/�t��jyb-FF{�c�5'j�?�?���ܭ��DG��Y���<�>[�=8����^A���b�Xt?1!�cH~���c�~���b�X�u��������z����f5�#�0dn�}���kw��6ݼ�)`�A��m�QX�=i�#5js�%a;���;|�Y�uk�a�b!�y$�R�X(ulԪ��uų��e.�δ�0	V�X��J�)�:s���"񗖥���f����\;�l��:y����^�ג��Ќ����P��1�X��7�cR���ʄ�b�>pz?�WV��I&1�Ȉr�rT�2�5��+�F������j����|1_(`鋐R�Ԫ�Ь�+vuv֫���"�T�Y�u����tj����Ĥ=
]�m۶��a2��=w��lݺ��ِ�ٳga�'8����$6�{��6�aN�ԆfS�Ua�@���BW�ha�B�T,)\q6�|vv��|ǘ���}d����af�HvC��-&��^�TE�k���hv���0���0�p�BGGG�C�����'�"tMaf����޾�����hjr�Rp��!~���٘gH[�ALm5f��"�Ʈ�Zqb�0Bک3/��i(�� 
��Q�1x�{�`p$;��' ��&�1tK\��VQ/�{��B\�.셽�����%�&Pg�7)�Xi�g�k��iJJeN��	��*K�) H"�Zd�g�j�d
�9�U)I *�H�� �*X�E�:T1���˳��#s�����������ɏ��O����/���cd�6�`^8}�#_.:��;wn޼����;<2:.�N�Wݷ�}����߹�@�١a:wai�����!��zݴ\H�X՝5�ת[Ɔ�mt;?�&� ��vdh���_|���?�W.�o6jV����Y^[�4��uy�������Sw���?}���ꫯ�A`1w�u�����ͯ~��[���ݚy��1Ԝ$�盾�-t`�l��h�Ԗ�����jՏk��u��΁<}���ƑL6F��JŻz�����~�pOW7TM�P�{�`����{��!UH�����5����l�m�_�v�p���a� djY� ~���iG������j(��/���Y�ۋj
�xⷌ���p���c�{7�T��s9)Pa)���f����,7SۨDLOO�1������u���3\U��?H$-R�)�B�0<<h�~CN��W�r���w���
B r�X,�����U%#��	}��''�����:���CѲk�JWw)���
�t`�ؕ�'�.8��M��ر�?a�>Eޓ/��_��~����ܹ��[wvvGb��u���ێl�+M���P{f��-m\n2�8ɺ`2T��������&J�Ҙ����f]�S4�0��-��:�Ϫ�{5��4֡�t@u�I�nz��x��_ig��git���R��ү�G,��Ho&��:���2Үw���u���ƾ��T/-�n�Ml�����s���2��g��ñ���\�LB[�ʷh�𓥥�*yMGꀼ�.h۲�UN?AN.�����Z�R,t2�S���VX��&S��_8ua����g�]�
s7N���N�b��G�v��Qb`��Œ燷oݾ~����J�6;/����xq�4\8_�Ŵ� R�<�'��Ec�:���������֛�piqud`��tb 9'�B��⠙4� 1ȗ�RGy���##�*'7�ꪸ�y�c����ͮ�ϑ����S"E9j�~`�JZڂ0j��<v�ձ�+���ӷ?<;����s�k9;������~�V�9uM�&Aha�f�Z�t���	WH$Z��独vn9��{jX�Y�tYYV+�˄�_�(7�feCH�Ń�ie��d��8��U,�N��^����"��4��ȓ�%�����Z����0#CӶ���|�~8��V��L�+<6l)�2�e�F���T)İ����v�����Ç��{��J+�|�T���T���?�"{]͒.�gЏ�?��:�C�&k� �n��+�+�0�A�F9~��}��c�e�o�>X�t�=9���7��
��ڹs'�<p�z�/�5�( � ����Ǚ�\[�tU2���r��>�N����������`�Ӳ�uyB\���֭[�(�"�?�8t�zQ3�ٳ'��!ƀ�r�<h\E��g`�N�-l&�G�䕵�.{P���hq����;�-���XS���<3\���,Ƥmٲ���*C:����00k�!��~��6��M�������Ʃ.]�D �T͹[��0�ع���d@�1�cؖ�1��=p��Rl��#!/���9l�dHv�q]�^\��;�m�i��,#��X7�B�@bM��@�[�Zu�ʾ��bة�
f$�m�����@��X�Y�L�ޞ����[��{RNxk^�6< �b�^H�ra`xHյY	�GG�?���O��]�̻+�Q=vr������;��ZD����A3�*�̜?~iiE�o	�{gg��W_��z�go�H,���^&s)��(���G���s��?��?�����P�Q]�6/�~���s�ĉ���o���:�_|��i�D�#�d�R�K���*;���L��oŏ�ٜ-)�.�o߾����B�O���`��F�6Sm" R�_�����Px��S�d�%��.����b	O8]��E��u��GA������ԑo��[:r�H_�ۍ��[]Y`�nA3���=�不/P�a\��>�*}�7tⱦJkØV�
�}HLg��0�#[��>�����qU�U�u1�!mαr i�T�J�3b	�U�D|m:8��ug6�o��i�>4�
	 tM�
Σz��|�L5���;XX����=v��@��F�x�-:�����$�m:�_����k<16��C�M���M-��ܤ4����ರ����*/~�h fH����Y��L�=q�"���XE�o3{�l�t/��e*�I��~vn�r:�D�O�q����	6u�1��DA:d��@h;>�@���q�t��tόM�}-���/�����Bb/s�������Z��QV5�#=Y���<`�+�V��,O�B�����1�m�0������`F�N&�@�2���F�ne�@.�]�^���k߸9��Ͽ���c?t���+	��Z�����F��� %�&&R�y� H�l@dş�*����g���E�R$���V־��CL����W��U��C�ّ�hx���KKf�,[ª�y!�o�I�a���jh���Ս�Ş��g�y�1�H�V���s��p �͡���5�'�iern��dg���.-��'�������\��4�� pq�ܘ��,cU�+R�i9�H���!�vےO&�6"ܒPK�	;�
}(�M
,KqW��T3l��J�#q��ҝ0��6���' ��uhK�XU�<ޖ��
l�bb�P�3;�\�8u�������+&U�lT�U032dcV�W�x.-���S�~����`��r���V�&�׼�/����nki�c�0���Dw� �IS��0�/���	���@�{ i��EhV�|�$�?4lwV������De	�%>�I��k�K�n���kz�4�}]8�a�P�,`��7ƈ�#}o8����R���q#Pi��k�p���z�``'&&n޼y����k��@�%`�0�&8�ĉ8 �{��g�Y�ibfp���I;u����@�딅qX��L�:�	��h��u��U|;3���1�3�w�^�
�ƩY�<����a��[L�i,]œ��@V���:&Ake��
�Ig'��fb��>�\��>7�������~O�:�|饗��0B���ׯ�'���%��
k#��X�x8��g�c�����auΉ�pe���R��P=z�t�V��pmSq@k�D�Ah�NAr��'��O���c;���� �����=�ۿ<7�W���'����ʺ���]���v��ȏ�����K���fs���]�����J]׮^��/-���9�s}�y{ff���3���ְ�U��N@XoH��ٞ�a&(B�ܽ+.R<P,6���Y,d\;��c�/�,�Z�s����
�>��z�@��}��ޱ��W��z&�a���-�@&X3���^���KC�c���������C�ÿ�����{n�Ϊ�H�Z�n%f�h+31h'i���Ύju#���b�f�Z�uv�j��zi*���"eY`��^�Q��粙l��Ļ�/q�^�_���8��k��+o��6྽^|��b/g����v����F1�vt�AJ�=��ֱ��D��],���W��F[V���I�2��g6K���	-���� �i��/�Ò�i0�`.*֣J�f��'f4�)�u�;��
1!C���\ou���s�(6�4���۳*�V/�u��c��C�O��r�
�
Lǥ�W�5��$���GAsQ%=�䓘�d�`}v9�u�.2a���}Y	9l���d�!r�]���jL�;�#d��i��li@i	���ȉ�D`JY����8�2ȷ��s4x#z!:�KE��<+:�{�i ��?���t:��g�=�=��i�;�k�FEgWWGg7� �
��^�َ�Q,����`O��~.eA�JEIM���0������E�������f����{�}l�ˉ�����Ȯ�;'��R�����x���>����>��de}�_߀F��@G�����~����zEY ���K��Z��8i�֖�R��*J�J��]��ԥ�Z�k�<�]..���Ve�
qa&�W�c�E���I.��l�'�Od�@�}/<}�ܥ+sI��%�w�g�n����e����_�2��Y��?�=�8"�`�˺,�|6�
M�K�̺� O/��Nd�A}}e�n��4s����G& {8��n�~"`��a�Ʊ�Ɠ��e��n�X���	_���2e�$��Lu�IT��a�-�!��o���%C���M��������J�q���?c_5��mh| غRZ
�#Sa�v�qEmd>sm������	��5ʌPE��6��!ZD'>T]d��s;vL{���Reay����f�5֚ב/�`����K߿���h�ؚ{�U���%{#���=���?J��
�.�s�����09
��l�0 � V�Н�?x�'��a���7�����_�sH|���9tP1�BwCҁ/�/�SĄ.]�D��1����P�p�7�qJM��s����W���
9��?~�(�w�M@S8 cƅ�wtt��T �ϺOiA�n��yra���/N�����ȑ#����4�Ş��1�5|����l��L8-D�ϐ~���3�<�q�̘@&j�p�`�o��o0]xv����~�{��zQ��J����,�(�)��"+T>�vɋ/���O<qr߾}�����X83��Đ��1H��#�T�'�S�����ӧO�0τ�M$ɡ�Bu�3�U��q>Q����ݐ�͌���y �18؟q�FK�h�v�;Vl%~h�A$���\�VΜ��(��{���PK�ʽ����ީs��z�XO����B>#YX�s�O��FC=�ʅ���[7��<�|���ضu}}����O�K�4����J�����}[~�w�����������7�	ed�����z��Q��d�����	\�����x��3�NҎۺ�fiU�ydw�vu���ƷM~�Ko�Q�ܙ�J����$��l���o*�VOA<�j�qQ��;t�>�]+Rd(q٢���d�C9oI�is-5QN�Z�`y0.��t&��VZ���=�������0�Z�Z�:t�����+[��Kr�|�P�d�r�\�tLj%lN6��|��w�������w3		ue�Z2�l���kU�#}@l	�Ǒ���!I)��M�!F��OQp/lbSt7+.|����\�vM��_O5�*���U�mE߄&S5���2gϞ���aa�վ��	���fJ�������4�)O�:�Qa�ir����.�b/�[,`�l�X[_ٵk�����󋳳w��*����V�,{hh��  yf�=z���Ɗ�������%��.�'�P�o���#����w� ���"u��R�n��tG8��%L���=�7���6��|�>j�wl^�j�V{����;�/S�+8*=<R>wY1Ϝ�Q(����*A,�Z*�<�\��-Ȋ3`�V6څ��̥�+�~e�mcێ�ccI��=�ao�6��o~��_��C�8�]Ʊ�+b�,,,A/ü��s��Z�X�1���}��cҬ��vj݊�H\�D�ɼ<�US�D1�;^M�^��W+@��d2��V6��qel/	}+N�Fπ�SnV*�ݢ���������w�(�;y����r.c��+��9/>�=��z���U��sS��k�>��Lb䗖�%5����k.U���t�5 �%�MXa�=!3"��n�t�OE0Pƞ5��ԭ���
�Z%��UҊ�$�DFHi��J^���oC 5	��H��������{����K�HP����3��04+4[�����g^���*��&���Vc3!ہ��R������D�*/�R-�v�)��@qF�:3�q}qe6孅�@��~��
�����wrxN���D��+��s�TY��0d)������l{��$3�'��`��<�4ga43a@��8L+Hڦ<�+�}�L�� kp6�z�q�����QJdS�hzk
;
MfU����͛��I��!���]�����<Hjo��#���u�������r��z
�����I+���_�*':��Fp��� D���ŷϮ]��C\�����ԯ�9� y;*]�lIA��OTg��͘@�����2�#E�Ꭹ�Tl߾�ҥK8?���b�d�Ή_2�	�\V�L������̼;j_�T>��o}7�3pG�ݻ��ŋW�^e%���1Ą�� pf���N�2��J��SJ�"s�S�LE�;��(����GO�A:�ϗ�b�����2qر�;Їqfs�F�ԬV"��(�M����։�8��\�rr����s++����읻����K}P�x�W�n%�cҕc����텝�+��ۇ�mޘ�-K70-r�`l�I�Ӆ��hnb�''w�)����F�v��A�H�z{s�����v�ڍFӇ���ѧ�Jy����9`!�;�{�"�7�����@+D@^ ���S'>��8��s�=��_�:��ߔ9<�P�yAQ�$��NMgC�$��2w��h#H&c��:����0[Dg���P�İ	�WV�ܝ�P;z6%��_�&�]g2��Ï�ڵ���ѯ~�W�~�Iܹ���Ն��]���`�c;�R�%��l�vF�._�p��?��-#�����a�܁Md�6����Ҧ�Tp��f�sy���V�J�\���L���V���2$;�Ot�O]u�r�)��X~L�e�3��3~><<�ݍ�pgb�ݫ�уXG�6U���y*)�J���j�N���!��}M��&��/S�f���5�^H9Ijhև��������o���Zmn~�Mu�	�e��4�暣ޔ�m�Nl�/}�K��{����!$$�=}:���:��3A�=��v�n�pRP�XH3�x&3�����WG��htb��Ԉ�}�1+�f�.����e�];����/���vt�D{�w�Pt�=q���v�K����K+��m�kb��GG���������w����:ӂL�?��=M���d́��u3n&Ţ�ur{qp��^+u�x�zh ��NN��5��E�Y�=�i!i� }��������}��GP��N�F��w&]gզ~5;�OcE*�˕������/}�ͯ��l@nKTm�6s{vaaQ�f3֛U�=,������Y�b�c`x��90ug^�l�\zbr[&S������~v`����F�yD���E*�a��AVZbbg�M1�C�o^#�=���.���D���!FB3�����a4�M�"*�#,�M��B�ݣ<6����|��:�a�i��4[kH�of�E�$��t�E<�^aq+�"�gwD�Fʁ��L$:j���M�����82T�1��N�r�	�l}��b�>9i�l����Ć]����B;��cU�=Xϙ�-��Z��
�l../]�ref��m|����z��B��)qa��E�&���6������OLa�Mz[�"��a�33��à��*�)XغssY��(.;������ �`΀�����Q���ø 	/	��Q�u ���0<��`�;��A�ٳ����)��{���`$RC���~饗T� �� B�Ԡ^��!��2:��-�$8N�V�+zI[�B�2�!a&ɠ��q��-fL�l�H�Јe ��&�"�2x����O<���={�%�cpڝ;w�$�$8r۶m�|R�؃���8ƌa���R���6�I8�I &�MI�:L����N�@�?9q�99p9"�(��q*Rh0E�� �q�@�z�I&���t�m��(�I��ȴ��P�%u������4�L�*m#e�I3����Խz#����l�Gb�tvwm���0���E6�}GO�K&�i>����禅���c)nά	���`���V�6 �I��mX�n�:u���c�t�W<��;z��5<�O>=qsz�'���ꎁ#�u<ʫ׮|��'�e�ٽ��+��?��r�������X��DQ�$0�	Gq;k�Y=2�-��Ξ���k��<�mr����Bѫ��:@�b?e�Y�F��=�:!���Xx���Ml��~�$��͕u�3
�ZzaGP3Y��{ާ�����"a�P���D������������� �.v߭�7��?�����_{��l���J*C��=RR`��Ֆ���ثKKw��M߸�p��c����D�L�L#ޜ�%�U���?5u����X(ْ�����e3��e�P@H:.u#ģl�A�뫫�0 L����VK�(�i�j6|�1���-
�0ª�N�̳�����SO=yu��)�O"�tW�4�y��{T]P�#�Ŏ�_ڄx�a\�z�1┮	�H�1BS:t�̙3���g�=�������942L�/|b:�)g�.�ei��Xi�l�r��R���j2��}�>����h'��lr�$:��
l���:�K�f�<r�AAҫE��Y�4�F��e���B#.)U�D<���@��{q���ʵk�$��kb�߿_�Uj�)y˙F����71>>2<:�;�V�*J��;v%������~�������������L��[�zjx���kXr�wo/���]�6����5�#��FM��g]���R>�U�hoo7�cp[cxXJ����n�� ��7+U�`���3�v97�E��=�R�򵙏��}��#�3,Wm��P��UaQu2��m��|���
�ĸuwɜ����\[/�|�81��^���*�z����|�s��P+�Op��m��c�I����a���m�%<à���c�2e#oy��I�T�*.�P�꼪X���؊�"f�����T�Z:dD��j7��I��qm�֢Ϧ��A�BX�(%�U�B���>����dwH2���7�<�}(I�>���ʉ3S-�����_n�f<Z犈]Z������+*�D�a>2Z��͛W2}�|OOA������o�6�V��U���Y&O%���4��N��6��& �{h��ή���:�dߺu+-xz�tz�+�?R�I ��z�a|��'�`
��F �(j��4==��$h�p2��z�k�IS4�b�v�*���P6�Z��ܹs0��oߎ���fN�1��8#4��~F���=�Y��%��  p	v�'��x�����1y�md���ڔ�v�ɇ��iB'��56�>�,����J���#�{�W��#?>>����O�Ix�嗏=���$�"�����孷�¼��[1?��������Iht�,����àm�a��k���;�1��t6NH���y��L�S�?���r������u��t�+�@M�Ƒ�;�g\���Y�\�����oL�wg�;�ȇ&�}�V��Ă��� %KA8Mc�ҕ���϶n�x	̜������\q`h���v�<ug�.~�HI�[�7�J��� �õ�ғյ�7+؈�]۴I��Z��0�xp0�X����Yv�����}����baey��T�69962���b˾u�����]c�v
#���˾��϶�n�;e��v����*3�o泹�O?�;<���f��j�:T���0�J���R���aD����>�&ㅅ�|.S(�:;�gΞ~������(B���6��A��T���ds�؏0?���>z{Psc�Ӝ��	è-C,�X0��vô����T���fnߚܱ�4ww�P�vv��a�剬���lT6`�ڎ��ݻ�kQʧ���u�o��I,	rV"7���nN߈ms��C�����ٌ�������nh`����L�ִ����^_�(���6���&ǳ6gu�N��(���05�90ؿ��6�a'O~
i)���E��]�t�Bw�ޔ��F��"Xs"�/x�������-�Ɔ&Ϩ�~���K��Y.�}�(�bi~!1��m�xP6��U��
{��0<<�o�>���'O���j�@�bVٸ	Bh�?�t�������}i7UC� ^����I�;��5�	��\L#�F��6q���n� Ү�tϺ4������/ M@����&�Ɔ��'���7oM�F��$���78`��0Ep�Z	o��b�J��>9�e[_���r�:;��M�]}P.�O��ccB�����"�����I6�e�3n�9{�go�����*,�|�ɸ��L�;~-��RU�EQï��JT.h�������B*2��$i�n�:���r���ΘF$E���;T,�/_�������T��W,fsR���9GQ�%���I)��޾gW#�ff7*�mօ�t�L����eK�z��ܝ��Ca��9�y$jUyJ�=C�%��*Z�Z�8^��mӮ�.�ٍՍ��Օ��!�q-�ު��#Yeг�x"n�,PE^+��)��V�d�S���ʚk��$L��N�:-r[X�$l���͵J'h�D��� ;d�V�1$i!H2��Uֻ�oUM�԰�D�D��ɭ�PU�N��W@��n�RӴ̝$�Z�H���q�5}iA)��$�1�Gp.4|O�J�3{�P*�A��DVrEa5hx�JE�X6%��`���5ً.�P��3l�� =�{|NQ�$x�3���W����ԋ�	T$T�$��=j ������C�:3�m�<������ZP8sgYß�1��6��T��|g|��q8-�L��C���ꥩ�Ο?�Ǝ���
��`�r�}a���8.H�m�+��`^�y��6�$������l\�Z
����`L;� f���KЩ�l����^;��%"F������7|��qfb`��555E^#���H�F�{��Ƽ}�+_���޽{�� �$�I�3�>��k&0�W��� q�s<2\�>|
���I'��>!8�ʄ��O�Օ+WX"�{d"'0�J��:Jո)�O����
��is`[�*�}�Y��~nyq����5�Y;R�@Vu�V& ��S������v�u�f\��g�3Y_YwmG��¼\�a���z�����؀�sr��n����A9R/--llT���[�Ff&*#:������_ǳ��O~*%�ʤ���6j������Zcn�v��8�mk��K��a�\\�;������ |J9������6H���X,~$��X�T�Fmuu�ҕk�;��#[!��׮\x
u�s�}�\s��D�b;�/6�U\Kſt����Sk������f����*� O���:���&Q(�F��������_|�e�5MJ�`j��c�����U](:�Ο���233w�깱�C��y,i�cy.�/��T.`!�q�U� �w���Fe�0m�X>M-rMS&�)ߪ���=����3������+�-�	� U"��X�A�K����RW�>���]�O��?�ٳO�1	��qS��A���zo ]� `��8#�%*]occc���gϞ:u�Nk��T��R��Û��M�����������H����/.c�4*��Pe��
2�R���מ];��V���%�ө{��.�$�'�s�������8q��G}�3�_��?�OL/g����O�Ul�#Bz̚{�=�p*f�k�{N�3�Je㽦�m��3��G����߬��;jG��t։>8N��w���|�g���X��<t���:�_��nMc�������֭[;:�O�������a��K�	�
g��(EWM�ۭ�R�HJ�6������tsf�P�ҿB��?�Wr����/�����;��0����)a�^__]�U�~H�ֶ�,���y�W����ڟ����|�ɡ�ݺ�J0�䟁�\�x����Q�u��+ K��r�w���M��2a�v�����EQ(���T������|*�|y``�k,�����}�(��<;�;�9�y�FHJzl�����İ�-'��AƆ&��(Ӑ�NA����bK8��5�n�u��D��gƄ]�#.
 '�R#�:����j�U�"�"�����6U;�u�3�.4GZ-�>������ �2ć��p&����E��-!�O��VP#��1Bz���F�ͬ�����QkVb�p�`���M���#K��U?�Du,zM��W�9vO��|Qѽ9�-ߙ_�ݨ6�z�C�mƑ���2y�&�Q�)L$E�T�i�;��X������IZ}��yZ�X�[�����陻�~de�Y���0RIh�!��rnK]�K����d3��T%�È�$��P���t�	i��	�c1.�]�tY��)O�gڬ�b,u�bfe3h++/u��ʊ#-�y/����9x������@)��4e7lk���d9�,=����8<?$&K�!�����:&���W�Y�~��-�ر��_�2�f�~�v���7��س��3�E��z_\�����?��O诽z�*��F�.���*L��Y������n�e�$8�U�����s�#��b��Н���Cų&�nPeo{���WL�$��L���7��;��c�<�h���qdd� Yp΋/j�K�:0�J�1�y���P{�PlW]���`����%ѧRlΕ���SK6��{Ab����(�02,؟� \�,Y�R�(�I��4d-�:�ߞ��yOoו�ӎ���b'�\�=h�l[�`����R�aT:��*���@(��<��y���cU�UV�6gr���{�$Z�;�&�ԍk���xll�op⳺��hx�B�S�Q����.T�ֺ;:W��n��T���T�Qȝ�p��S�������?0�;4�z�˿���sk�-�̶M���n,>Dn�$j؉I� by�������X8w�`y�D��.*H�C|;��M"qva��o����3X���)�xiQ��5I]�*���6����,�ק����/,���1�����ΫW�OMMѢ���y��Kؘ����֍�kkP���}�f҂!1�)�d��	iwL��t/�((����^�i��;o��k�۶O�ڵ����Z�ͺ��'^� �d�
 �G>���?�'��RY߶m;�Sk�{MA�nj̜R��{�w�<�z�(B�|�w�\t�g�k3�Bs�b\������^�3�"��!M�M�SXu�����PT�v���a�І�:'#���%[fue�1�t��ކ���ӛ�s���b�A��ka*�a�i��~���F�^%�n��a'�G�}��w��!�5m9�u�/���(�H^Gh�4�<�<X�x����#Ϊ�"�=VG���[ugs=����б�v��6�a`^ñ���C.lG+o;rS9�������=�=��"�������tG��Rl6�s6c'�q�MM��mf2Y��K�E�^BW��yTE\�����\o�.uK�L��3������,'(ި(���zZ_Z�,�6��;�G� Z�KH�SQmZy��P�N���J�"&�@)!�i(N���c��..ͯ���I��.�1�=;?hblU�Ɩ�T�����.�lJ_Z�-^������`�4΂ĹB����6�Y��L.��ϑ��Y��z���%�������fGZI�ʁ��I�n�I���P-_��B��fK�RA��D�%U�O��F����6�D�iyhfm"cz��ő��7Or�[!�@�v���dI�Z$��z��^�T�"4"�v;:�FS4��Kn��0��)�gy1���#�S�Ts���滺r�� ��OQ�%���mc����Jo1+��~,͉��7�l�;}�RDF�f��4ӌ����5�������� �U0��+�I�Ad�V,c5l���R�w��D�9�<�2#�ׯ_�OpZ6�Z-�7C���N2�������)���6$L���9�#�uE�lR��agO�u�� 7oބ�ڵk?.!��/�Zr �/~{�pm�<8 �)�EJRp0�g�}��g���X
����؏'< �+^,=�����\G���ك��y���S���I��޷���.ee���:���a1��#�!Q
�dJz1�͵�!����̭b�&��Z\�[c o��&.w��	�:v��4{��G�2�'��r��΃y�M��}�y˺��z��|L����h�Ǵ�s�14�Ǖ��Ƒ��f�WdŌ-�t�)6��-D?Ql�Vw_/���H������%Ծ��y��/"E%tO��`�E�qjb	D��~�i�10�Tw���x?:2�?�����W_J�����?��?���k��Z�v���������jX�Wir��'��u	�Z�[���?~�;���@�Я��o�܉!���bq�r�F���?�MuSj��jл5�����<�k`�|��_��&���u��@�as��mő�oϲ3sk�6V#�<��sXQ���#^:���<f���C�6��e�S)`�B�Ƒɂ=�L���X^\�p�sg�Ww26P�՛����˜.���#y��ݻ�������ɧ�8�o_�!�6|�V��|����\��Q��(a� ��^0!�@F2�S11����S_;�5_C���į0{��)�p��t�h(B���p�&ȱ	f�(⳿t�M'�5N:EY#�v!��N�2�_N_Ӑ��n��Zk��>��8��.�c;l+}{ng@�lHZ�X�:�Ѧ�����xG��@���kQ6-r\�!�V&}L�2ib]Ʀ�*�]iq<HǻN�@���x�Mt�̺g�	����SmDa22�%�+���vuwת�P�8�Ϥ�b։٦R����4�A�'��B�zw~Vw5M�P/'�_q�C�դ��BX2�}��%1u�c�)I��8ye�ɴ"�i^>M�<W���1�	��b�2I�#dc���Z�C�0C�9��f���Uo�P*���b���0��_�:[�<D�Q��\I] PP�sjU���,��D	�	"K;����o����@���=�����+�SX�al�D�kg��V�gpe��ݬd	L!�SE�+;}[%��r1]	���P[���~h�9^�e�%���&;>�V���P��7��<i=f�Ǆ�NI1��d�I��A[i�@AB�n��oP6��W�֢�W�3�.i"2�
<��<0Q9�`Չ��
\C�_X�"�t���QѦ�$��7דO>Y,d��[�"�Z������Z�@>[�= ���3I�̦; ��d���`�S.� Ɠ~f����C�e��Z�
ZdC�2�V�&�6T�n�Lpr����&>� XwH.��0�)���r#���9��0����!1�'�|�
�v%a���/^�Ea���,D؆�՝� 59f��r����N299I����Z2F`�p�mqBՂ]H._����n89�L\��N�U-�ۙ3g0E;w�Ĕj`������z�2o^�c��"����%�8��|�lA��Jn@�q��,�b�p��^�#�C����<8\�^x�'�]��{�$�m~�_�I�}D�c�|�+�C���9y��J jq�N�5��2n��U]E�5C�G�]f�SD}hš�mOgBK�!��.C)x4���t�dFX\�|F�r{=H�����tjR3iPAFDmz�J����2f(�T*�xZ2?�8�u��^޲�ҙS�����o�Խ����7���ߨo�WT�GF\:�d�����&t�--eMX�Պ�q-/.��⊯�ʫSW�a�cf~��������=&�q�ğ�}`���QSCQ3�s�0d,�T�  ���Ɠr�jy��q�˗�B,0�;s�&�#�a�A0�W 3�)\���6\��ͽ�:�"�����bsa1_���4$��y��S�駟b�c;sYbSӰ#C3��)���msag�v6�Q�l�8������ݵ{��7����[,�?9~B����\ԫ��UT����q`ee��~�K_������i&R�및n��5�=�i��bjd���m^AK����ɔ�����6U"=�^��m�%��)aS�2J�-��YߘƺZ����>c8�5]m�w�-�QF�A4�Q�'�5�i�4��z0�C,3[5��Ca�f�.f��jB�t�h�V�����7H�3,��hQ�tb���(4K�e�ͺ�_�{��t�B���'���f{��B��h6��Y�eqP;�N��w1�CE�AE�c�*TWL��H��X�B�Z����5�5縞��p[�|R��;��
4rH�{Pń�j�+�o
��e��-f�Cc���A^8M�G��(���q��{SM�Y�OUflrJәV�����NC�S4�*� qn����*���X�4,E
���{{:��<0�?ْ�\i������p�;:r�Ѐ�M;4�0dA�vݭ�����{^s���]z�r��xC��U�(F	�"�M�b���A3n��1;춛$JB��*��XȊ�A��;R��u��lC�1���p��W���H"�~Ö6D+���n!V�+�+�7�O_�0s{fm#�BJ����KT�Xq&D�<�'�3���&o��ݳQm���*_��v5����%��Rd�/���Zymuqqy	�]ΐ_2J�̎��ݎ;�?��^Yw��J�]kh'�B�$rd:<� ��U��ţ�������,`;��x|T����e>�IJ�P��ҩ����H�C���lf���N_�|�ƍ,��I6�#�w����¤����:y�$�yꩧpE����Nz� �T�$�ɘ����oM�BVk����G�v����޻w�z�[\�w���ŗ�283p��qVۃ2p�A��v����q�!;њ��$��.Fs�PgƷtM�J
�Ð�?C�Ҹ�T"��M�R��묎`:&�F'k��s[�~)�o�,��^y�W_}s�	����~�m�r��Zb�[</�P�ΦĀA�5ݨ:�$���;b�R��l]\���5o�Ts+��r�6⽬K�N��7!#	�GB�o�.1]�������������K��E�,xɵ�䪡�ivc�{|�y8t�>Ě��Y��Rww�p��0�������gy~����w~���?�80�ze��T\Y��r
��KA��n��c��������J�R�<�4�3�<�؟��'��g^z��l&�-CK��H)�χ���4�FG��DH�U����a3�x����Ç+���b�P,]�F��'�xZl�ȿz�26#[��BA=��b*縅��0�E�� ��g���թΎ��r�i����۱{7��~�%�3c��J��Ȱ��_���ϱ�¡��toI�yr�Bb���}����־!i$�����T�a��0���qsff;�#O�Ʃ�'Ϟ=k�lC�ƅ�o�~��U2��^��M0.ABm��K��i@��
�2��+\���Z)mI�-�+p9�{}{�75�����'���n��hI��GUmH������Ԝ��ix�2`�Ò��HgF1 @��P��r�C��Od��j����ω��c�YP�&,�	��Ou/ �I翥i�k���蛞o���&D���I��Cl���e7}/���粅Z��V<==}b�nFy+0�$� ��^��P�1�n�J�ާ�N�6�z�ی�<?��"�C���3�M��s��kpb��-rY���\�V��R^Z3�"�,��1�PB=x�|ϐ*Y��>(X$�I���D�b� .c[��s������OM/����@ǗLE��,)�s���!�|�6_\:�o+��L6�ci���J e;h��Bρ'F�=��,�ule;���rkH�����]�\������-pU=�s1s�M_,�8$��8Y+#=B��61-X��l(��K�J�c�L-�͐%�m1[.����51U;`�ĵzՑV��R�r�Zmtmy������ٱ�Ϗ���	�j8d�#��+i��Ju��֬��U����&�����G�MV�%���t9A�����*��ŋ�lib�x�h���y�9�6i)�M�`!�t�W5'��F�V&�H`�a�АŞ���81�������=Nt�Tr����^�v�tzQ��$�Q��]�"2)�`�f �M�0p	�4�6ݟ���c�-��4ݨ1M� P�����Y����!�;�F�j�_P	�J0��O0��*q?�j'���'1�+W��{,��	K�T椑S��R��d��m�����Xʜ:�20���b����C��e`D2y���
�70�h��;v�������}�t���vϞ=�I�?�#�aN��#1�^P��6p�[o�����8?�d?%\����*��}�����)`���mر|��q\l�>�ܔ���3�3VALRO���e�Hoeۆ���$0?1��Eċe@.(6U��\�^��Woq���[H�}�Sě��M�J�ͺ˻6h�!�.�F�J��P���u~���k�H�z�����b�0{{��Ե�۷Yn6c�=}xBãX�9n&�9�cz%��M�q;J��wU`�r	{��l�(�lı{��ju����ˀ��OA�ُBq��2��\&�eO?.Nu�ܹ7n�Na$`m�)s5�nU/\���O>C,("L���<�h%�X�����rH\]i
,�D�g�����2���ٻ
�K!֯�������3�vI��^|~��%�����ڹs'��F�`װ�#M4��-��.��$�hw21	65�y���։�'������z�b>�˸7�Marp �v��wg/_�
KQ���2 E�i�
Ӣ�l��j`�c��Ϩ
9E���2�:�aYjssq�2��9���)m7?Hu�>�?�X�S�4
���h0�{*<M��C�>���o���
i;EPK&�E�(���
C	����b΋F��g&�0ˎ�:��u�&J�	s���F��j6፴�Ϩ�&>�M$:�PO݃�����?����j�����箜�u�U�Ǎōn3���FB�(f�H�&:�ǬNo�F��$���U�tt�>\S���"d�����M[Y-�D<Ȯ�ؼV�2�dᅪ$Ȓ�3v�5T�`�M<��X%K�X5C�i��iI�I��M�NMb�6AQ�RM��"��f����l�v�sN���aD�i4ubîس{_��������j���8r���C�EbY�>=�B�h�7I�#泹l&�B;F��:�u �Z1t��lT���X3�0�u�yy!�x;�"C�tT��q�K
bTH%r,�Z#�m(�ͺ_����2��F�`a�+��I컹�"����a�	C�^̈�!$=R�$�$���C�E7Wפ+B$y�,�@�^L7m� l����6�]�g����y���jU<�C��Nc�/����p$��u�sXN���;�`�O1�	�$�%�V;��&�-����ƚ�aa��JB�VW���J"����s���P��nl\H��j����hVR�3�C��|\��#�^�}wwc�)�P�S*NȔY��Y��d-�k766F-��A8����8G��4�E;2Y�O�D)L�Cf$�$���r�O��a�Cx�% W`+c��1�����A���h���p�8o���r�6Z�,&����~�)��o)"_z�˗/ �߿�k�ݻh�F��iY�
ly��Q1t��`"3R���HFWEĥq;b2�6.���3���$��/���0-�@|�Ko߾�5K0F�,>��c�����<x�|:���X��uB���V�B�����8�O<A�@#�//)Xp��|jj�i�������A�r��S�*\W��AhF,M�cX	�D����!���N�,��cwm��$�*�&�: ���:6?�FƱs���+z�>G�kŊ��4���y�)Ce��MU
	զb��v�𦶍	�7�TKV
���.��j���t	�BolT���������{��'��3����hy��F`D��Ј:��/��=BƁ 4�?F�{a6#�%V(�:�:[�ƱTF������'N��;� ��	��V��o���q_�`��fg����M�?}�za͈XS�bGŖ-zL`��zO���x�ufI�����(��X�K�Ѿ}�P.�+l�X5�a$�)X�����+@Μ9Ў�7�T�I��\�W$#i�Q���\ߨ�8��c�ݝ_�1��/~���+�	��5=�-��9{gfc�<62�e|+f�ĩ�.\:p�@oo7𘞧��9�`d��̍�	�'~�����=��dX&�1&�S�8T* mt]ՖN���zڄH�i�9�7�����v�W�y�]H��-[�߰5Hܟ�Eh6�_��� �zzH������!h`���MHJ���f{wS�x��6vfrv.�����x���Ҁ�$V�j�#T:�6.�a�t%��G��i��i�@}_�\Ϙ�TZojA����6�A�1Ϧ ��J��8v��/[n!��sd��:�"f|���5�'a�f2I{�1��U�\k�P_�/�,�R�R����"%�4V�tG�M���rt����A��ڱD���#[$���.f�Nk*>2(�C<8la�xbk)�+��\6��T�Rob�1@��%�4�8�:v�ȑ�ѱv?�DU
53ۢ$�a�AX+��;w�����$vG͋��guQ3�%%Z)�i}y�4���@,����� .�iK�)��pm�ndY���4k�9�c�ֺ��(�j��c_z�B�a�ì��B6�:Ҝ��lM_ȯc�	h��41"'c����cΊ���FP���6��Ᏼ�S����\��V7�zЀ�5��X� �] 5+/���6��5/�&}��g��������S�a=�X����˽�>ĺ�L�����+����E-��[���g� ��oM��K��%4]�6+��!��r�X�QS��P`���E��������F��Oػ�_��,��H �a�l۶�$�̗��¶�x��s��+egn�-Z?d�፰�20�mR�2�!n��NM���8L���f�>�"�	�ˆ^fFi*Rv���v��pBYF�`�H	6�x��0W���`�`.�={�СC�Q����6l#  ����� ��sf	�W�w&�&����s�=�',3�C���D#�[`0,q�ɬM�{�r�p6�U-06@����v����1Ӛ��@_���į��9u��Z9�4��SD����P
�3�`���Ü|���>y��w���g0��/��2&
 ��u�",9���%%:��[�3�S҉��'F���������H�Z���bڭ�!g�`� ��'�h|��mۀM��JWWW�JصT�$���2RA�M�V���~t���!PF���b���~�����;&�Cߜ�V�YAA'�NC��VP*�qO44��P�u�++yrB�Y*
���$�Ե��je}����$��W
��޾3�|�G����Lm�i��g=77GJ}��+0���a���S.�V��a���=��̰[q/�)t�n��	qq��E`!���[�$C��( ����1�8^��c#���`z~��?�)�`c>���l��z����7�oNNN¢�*�����M�6�2��*���YZٸ5s{eu����}��jMQ;�bs�%����Ύ2�>����w�.^�7>1166�V�i��NȂr��z��M�;ab�Cֱ-���a�	g� ��8 ���lV����CS�t���k\���IV���^{�l���eJ� �7u}
�Dg�6�۫���4800:2���4}���=�S�S%qH9Lt}��eHlz1��az�^�J��o~���=�t�&��Z�t����DW�l
am"�O�tu�e�`�v��2!M���b�(��u���ɨ��
�G͋/;����D�X�.��ql�6V���aߋrT�Sw�����0#�==�Vb��U�u�qTC��@�����d���-T)� ������rU�SU���ܚ'��"9���|Dc	R��`�V�ie�Hj@��I �`�$F���8DyH �U.�k�Q�m��W^y%�#���T�Q3�X[��$[,C5�
�ޞ�B�(N�8��{7�����Ptuv�:�4M����!�Ws�METf0;_*�J"`�ROO�V-�U[k�:�r��T�%�i�.�l����ͅA���3��
4s M%	������4!�
9����cl`�}[U2Ko"�R�0*��fF�㊅�*CKt�!���dl3��.�0|�X������R���$Ul�7������c{�?}��R��nG8�Lr���5B��+�'�4]��1T�Cgu��l��Ԍ���Ͻzq��\�|0��zSg�he�� H��2��Bg�Y iPA�55I�iN�X��	��UM�5rDB�ㇰ'p �XX*0��P�Q�/�t�q��&�qZ`s�ĸ^��&ƣ���u<��#
G\���a~93�?�j��.=\����߿?�����R+�����}��8l��}���a��'H��Y�P2�ᢘ�cǎ��⋀ΰfV�"��o1Q���_�N�����#G��E�. �.f��IDL �ypG l�?�<mt��½c����F6&�B��`?Y�3��}��G�.]"e� :;u��Χ����1۰Z�O���8!�!����|����}��{�c9�&fe��E�1�HI��K#���V��n.*G,����I��ff�1u@�ݝe��%	���C�)��"'R!�d?� �fU)��y~������`�ʡ�/����m�YM��I[�����w�=͊�[2�۹k��={���ޮ����t4�5�UH��B6c+(�#L0B�Mɟ��N�B�
N��W�v�z~�9��/{R�P��Ǉ <��VnN��o��Y3iuZ3t�p�Ī Qx������~�������c�'C&CJ�讫��)���f���E����G?����=���5��CMm�m�[��[��a�����_��}�N�>���N�4t�Vzꩧ�φ�ϟ?Ղ�}�ߊX��
�t�R%m_Z�NM�e���L���L����~�α0�'���n݊M��DN�={����j�q/]�8;;7ww����'�z�����/��u�.#�'%焙��h���~���0�q�x��bTx.o��&�o��o5�"�l�ά+�4�r��8�qt�({Q<��@H��D-��y�ƞ3鼬M٧���CcP��Zd'J���C�=��3�Ο��9ú�]r���M��!$�ɓ'�1[�)�p�'�*dG���{"�؈�[�n1 sK>X��{���&�����tiB)��A��t#='�8�.���r�T��$�S:ꛆ��	�}���ON�m�`����o���厞|>G����ǅ���v��=2:Dx�{�.��H>|��A(,�`���,,,2�P5�
ӄ%��L��-�!�-R�Q�3B�ӪOЋPu�1�?��4���:���߾�wϾ`03�H$$Ҥ$ӑ�e�������R�\Q�?�G�Cq�]��JT���+�l)�dk�I	BA��D�$�Y0kO��r�����9�s�o�̀R�/�<�s﷾�9�9�9�)�rM+���'�`��Fa�2�eK�d��4'KZ�+��)���8�2�i<p����Z�FBh���&9�s���k����17�Xz4ޯV�����[�۽|����ܨ�X�&��h�Rk��ܧG���m���Xddc�s���a`ݠ�ZY��*�pƷz{�8Y�Ԓt��ݹ�h��XK�x�%�������@��[RזQz�&a�i�ׂV��| T#xٖ������`5���֊Į%]s�8�����J����q*�oIN�U��f��8�T�RƤz6��jq?��e�(�h-4�=��Y5;��A��EPo�n����a�
�����X�#'�sg�uK�(�����	�O��a�<y���U���;�(FD�^<Ų;+n�2ߎ�,I�aR#I+yn�%��;�����|�Ã;�ٖG��W?�+U��ߥŅ����h�FK�$sc\1nd�=G�v�͜z��p�)\2��9̑�����aQ��x��௿�:�9�2sf8���
��������J��OLr�����ud^*�Q8`��?��s�d0_��dр�<U� ��Q�İ�2�r�e���W��U�"���"~O�Ŏ#���b��a� �c��X����8���p3$�o��8%��}�MF���d��w��? �!����{!%_��|��gq�8;~��	H�k@������P�%��w����)������~�i����0IH�AE2B&@>xn7��1B��&�)n���Q�/ҹr�����k�K׉�+�s��Yv�2o(��Tt`N���� W��lF�f�I�/��T� ��\~&J##4��c��w0�a�e��\�xena�XN�r�Ҝ8	q��SQ[�e,�!�/Ҋ!��s|.,�,1]��f���%Ȭј�,,��e)}X�f���Q86	�����.�����6�u�י�E؞i�F~�as��|�M3vVX����cG^���$��G��l`̱�����t7�tGF����Na�ό�h���P���®ɦ��T�,����:p8����������<�Du"�'k�^����>C�1i]/�t^� a#�_��:x��r����/,<���(������lZ�6?)�YXX�B�jG�����׾���ƿ��w+�j�3���l[��ԾYR�K�G����o4�^}���_;���(��������G�T�"���D	0�c�=��/\�t�t>����o������?>٤DZ[�>fS+��<�x��u�x<������k7q� �g�<�~�V�G��;q���������+_�
�秞z�����ys����N��<���Y�l��Z�^��^$��8��S o\���sK:�����{���h�������k؆¸6��ؕl�S`BG�M�� ��<��@K�/DQ�r�V.�3+����@)Q���I6pZ��ָ�E����W/ߺ��:��g��u��gJ�
t�^in�n5�^�V6h���~p�@������0�E9�H`xv�v�=�Q��_�Ƣ%w����(Ȏ>.�j�_��_#�����8~�?�w��b��0�A�i~���/�JdY�@�*R�����>�7P&��D��C��A|zl#�� �rg��K�yW�_�� bϲ�����?���>D�CB��W��[/��hԘ��C#�C�����c'�|��O|�� Do�����y�G���oɬˌ�/ ѱ���9��uL�f��[8���9�i���f<6c`� rY*�M�d#p���Zk̵q3�zm��B�Q�J�ys�R�]c��y6&�$�\���S����h2�΁�� �������_�g�Ӄ'N�X�w����(^XZ��j������8E<6�E���yU�l���}�V�!��Ӗ�����C��q��I��깿j���x͹t�����c
+��������n�i��P2���.56�MD�c9�?�/!kԤ�C�-O���b{2,J�QT���d,�!|�Ԡi���!�+VX.�4�]��|L��چ|	��vu�빩�=����B���n� ,k56`I7��V�I/Z�c禣�r͈����|s�&ǐ��8��#��
���8T�-&JS�� �Q~�Z��|2�;��}y� �0p�[�����Z1������>�|i�0�c6�w'�!CZy0������Ώqf�Θ�gI�=�,%�|�'�!�y��K�����
�@L�#��U�,dUi	��4��	Q�~�mV~x@�δ���{����pL�0z5|�}_t	�0U�
�+NM��7E�=>��?Ʀ�W^y��7�d�Ż��H�
�����l��@Rd�����*T��򗿌�ォ�8�W)6�0�p�/}�K�H�+�� �Ɲ���U��?�cz2@��\D�|��(%�ގ�q {^O�W���hY�!LE ��㼸_�k"��\Nx�lJf��5L�y���$cY��`[�ü�'� ���JP[]Y�//^�p��5<���E���3N����7�Affe)zU �w̭����a�"�s�g3��Td>^���D���X|%<�]q�B2g]3.����n_(�?d��Or��p�9o����2^`�^�?>�[KBX�_�^��h���E�E��������@`�/��d$�ǎ��=�V�Z��F�{��������E$�д����_zD&X��`�׫��о�0���jڢ~T��LK�g>�7��?������m`�?��W�B��FHvm������_��\♜<y�G~�GN�~���S?�#?�����r`��Mj�Z���
�:6ϕJ�ŋ`;������K/�t`� �kqi��wD=�}�Õ�uK�6� A@��#*��@#�ba�8R3M\�*.�?�G�&�h��g>�c����8>|����M�жZ��%�~�H�������ob���@����|�O��Oz�s��A�hf�P�ʼ=K���+��^ZY��넣��͛0���TX�����d�;�y��^�mԖ̽)���q�i�%&� �㜈bv����prff%N�-�S����˕ɥ%�@��4�r��Q�.��q�b�:n^Ɯ3�3��r��~zk�t4��qd����u�������3A�&s�d��k����O&6���q��r}�/^"^4)�=>� ����8$Z���{�G�߾+3���8�sYl�e��@����5�EB��>�K
*�_�r����6*��>���@����������n���l�Jş�d�a O����<���R���(�(�g����[Q�񀂂؅i�2�@�J��%i�>,y8��f!���%��G�A�0�r�Е��k+v`��CTL���� `QQ�U���L�+1Fy��jc�(��|9����IhT�`���z ��hե��՝��8������ R�C�٪c�!�I��|�j�l���.�Ձ���ݳ+�F�ݿú��z�_\���\���K�j�-���e~[4@�0���Zm���p �ם${�[s��p<t��`U��*�Z�"�|��t֗����Td�;Y8��k��k���X�k.<s\?�x�����8N�x�5�<�N^t*���G�d}(f�p��h���$��6 PZ��)#���Û��d��P�ks�N��u��8�l?��������d�ǹ��
1�Į	�	i�7��4	�܉Ѵ���(8�%o%��Ȳo�ؚ�i�^xFcju΀������t�Y��"ZX����N�D��Q�i����4�R�X�H�_7�X�K�W?�͵,Y��\�g�	%Ac�)��fǲC����ܤD8��{!db�N���qP)�1�u��1@�8~�M��� ���
ķ�B��e��O��Yd�=�!�|�{�#�_A�
��+$8�I�K���dq�Z���qL.$��]��RU6g��d-�a6�+��A���Sz*�,8XgX�Ŀ��[)��>��o���q욡T�8�B���.2'0i��a6C�vwnn�������E���Z���74��;�Id��H�/Ѥ�dՍb��=U $��$N/��"�	`4v��R�j���dX�D� ����urx_������7����^�����F�$3�4��ت4#��>���"������gz�G~���7zA5+&��k��T��;��F��[���ApRT�4����k��8���{�{������8��7nn�����?���/\����eR�D��4��`Zh�r(�*�FqjDV�~�����¸x�>t���X�5�z��E�Qc����5۳��'�x+v4��^z��{������UCL�n����5�3Ɩ�W�g�O��O4��#G(bA�~���?>�i?�������ck���󯨵�ղ���=��?��?��G�CL˸���q������{�ѿ��?�a�ߺ�����V���Xn���<��c8�H쾇~����~��~�g~��y�s�(ܢ@w8���&z�iF�q�k�7/\x�^ �)
+�X�K��(���i-ß�?;7�#�H��H#Z��'s�I,�br��qI1���*]��#�Vُ�1 ��^�dPk�`y�j��߭�!"��td3)+++"�1J�&���~�������yX�J��JɠLa@<��ǎ���۲��49J�M��
�\Etd4�Jc+�3U|R�v��O
�,i����u^�6Ք��5i�Wό�"yY��,�]n)�z���>P ����ŋ��F�u���ޠφ[��X�]H5#�(S ��k�S4�Z��7��ʧ��۽~}�w�{�O��҄��f���c7�D;�I��Q3�Nn�z���<Tn���zF��=ɒ艇>�ȣ�˫76o]�r�V�W�woI[�Hd]p�iV:��o4k++X���[���1��y�y�F������ֿ�w���O}��W^�9e�2�h2@O�K�j��V���x��ܢyZ�����pl�!��C��Iaíʍ�ں�������"dF���p2� J�M��k;�>x����� !	�S�����Y|F�����@��c!I��:ޖ�s�9��5��8�� ���|4 ��;��W��4I�Q�u'I��ҙdK����c�Ѫ�*�N�bǸ�L����Xf.bdRS�?����PR�v�V���d��(U�\F�X!����w����ɒ�Ɨ��8�ey<JҨ�^��T��x2�k2z^�η-5.���4�i���q�.z1qܜoT=o����>Kތ U�S�p3����ey%�2�{P�mh��	0�����2a���0�!��+'
��d:�(3�El��!eɦ��)���F�`�LX-�.YI$1�����x6���R��ؤ�S����)I8>|!a�tp�"^63^����L�EA'�"�$�c�>5��o��9Q�0E���. �F��H@�?Vx�`�~�%e,U$$�!�l)����*�0� ��`-�3���p����U�u��J�QP]n�6L��'R�E?��,|��/$�1Ʋ�VWW�z/_��+��b��j�3�Qu�[�ؖ~��(�Z) ~<�ʊ�$jV+K����v��xǚڈzEҁ����ݮctL��F�1�c��`��A�۳$�Lb�,��p�kL���؏�*���/���>և��F�C���C �F}n�����QU^�#�x���T<�22O�-1GDF�-ܢg�b�8�W�k=���������
�k�},��Z�?�w@VP��R&6E��`8� z�������e{���}�s���#���B���N�8�G��}�k��ۿ�H���5�eitS�\��hL��0���ŕ+�~�� EP����C'O��U��^�8B@��?�����{��!�a��3�<"q��PI��Ȟ{��ׯ�l����wT���x/~㛯���X����b��O�E<�_��_��_�lU<l[�#G��c������ϳʍ���l:5��*��u�_��.�_qF�uׯ^�n[��d�t@��c���F͸�+�=��(��(�֑7;40�1jO��l��(+˫�vm��`i9�8���=���y�eϭ���[1S���|��@�~U�{���û`k~ef~X[�v�q�?��ﱳ��b
SO^���H�c�o�̭z��&E�|��ń@Lf�%����!�L����!���M�ѳkސ;EӦdO��i�Jm(�%-��T�����v����LF�=x������ŋϟ?O�:����y����z�ĉ�W�b;`�a��Aa�c;�;��>|�3�i�f�6��n�� D4.�3�sƛ�|�+m^�Y{uq�����O|�,�����������/^��"��4�Y�Sl���WV���${��0^$���ul�x<
|�]�����������sXW��k̻D�9.M�\�?����W[Z��$���(�� ��M>�(�$֛��0���q�`1�bSy|Q��q�[/�yry�ɳG���ۻIW�~�X~�U5^Jҫ�d��c�:���t�����ƜW�^#gkk����n`o�^G���C&?����b߲��%Q�j�w�
�:�X��2���p��0��G<�͸y>�SPk��w�Z���ԛ�7n�T��A&@��E�a��z#+�A]~�x26�F��m��Bl	b�6w�3����*�����^*c�dE
�֛1�pl
�A\e妡�E8�����>P����$��ڂ����TK�"ػ�2änF�g~h"U��<`Φ��+�&]���X[g�Fo[)�į(S�Gc�.������&�P��3�b�*��!��a�E�ͫ.���u�>�9TN��q��"лs�*;?X�����)�<���0)�D/_C/ʂ��4��Z$:�`|F<V&�3�~h>X�Y�����ݷ�,�0Hb�Ixx":���?�oj2�(#�L5�T\:��-O�ÀL��0�����骉��`^�KHW*_�	�j��;q$b)�f�� �Rލ��2�B��]3YB�!6\��ߪ�"hb&t;q��y�
�7nU��Z��8���՝l�e�p���S�;�2����0Dx�{ݝ�@H�~��|8=����E����[7�f�إ�^q�\{�ڵ+���'�o�Ϳ���w��np��>�ưJ�����O=��mmݴ����p|%5�;�[5A���֪�u��ǬJ��$�62���/]����wmnn����P|��C'��%����3�KC:}����DB E8���F�u떪��j<7J|A��k~뭷�`hP`V�����p�g4����wnl���_��7���IB�ɼ5��c��Vk���LY\ ��;	P��~�S �mɜ���q:i��˹����~w��f�^2T)O� ��j6��8�/��S�={��o��y2RE ���]�������j�v��By_������9���.^F���&bQPQ�i���[�㵳I�љ�l�6���=M4�M1�`*���,�
&�$kn����� ��َ�ja�;�6�:�шq��W�نC��TZ���:w�"ܯQ��ա�!UO7�H�8��� j��I��s{��W^�l3"��6���?~�8G ��+h�/������R0��e�k�V�!�N�jV�y�����eV�C��O}̠1�W��P�����o��~T��`<�ϰ�J��R���(�C�n����)׍��!��Pc��n������|>km�U�#4�c3ۤ�l��X�LʢQ2�Ʀ'Ա��l���=��Ӌ���ݧ����{����W�\k�[q�J;��l�D:�=y��*�қ��;���1��T����{K��7on��F�!�,�����љy�#`=IȺAa��H�Kq�?~p��^o��7�����x8t�����#�2(���|z>�"d
,.��F;#+�;ݗ��j>\�Ĺ#G�jU��sG�n��Iի7�)���;J�p����Tٳ^�ԭ�"�=vg8(��w�V�Z}1w<�%x�Z�S�w�v��b�J�ʆn�/����N���$҂����M����`,Cʁd�gI�?��kE?t���%�onş�t�Ud^<޿�>�x��I�v�V�gi�7�g��'i�i��.S��
�q�d���cԬ<�x��8�U/��ʔk]#W��Av'�-d^�n�Oa�$v7���"
K�tZ, �>Ay��=g~�Iqe ���hЩ��<=3Iڸ��FC���j����&<(��Mt;��� �`@AceU��u���L�r/��V�� P_��X��50}[����ۍ�*���Z��Y�*�ć���	'K�x�,�P7�R��8Ʃ��G`9�d9�G\�
Iz|$���o>=���H@��C$���EhD��B����w��Qh�Ȑ���a3 .W)��o�20�Xi���f�A s$��w��f�F�I����cIl�i�q8l��ÇVV�;�.�G��I�X��Q��Yx��������p�����o5��ppV���^�+X^Yb�6긬���q<��v�`uu�����8 �kׯ�5���N��� !���?�o�z�ĉc'O���;Ｗ���S��o��܅��'j<��#2/�a�����L��¾�H��^o������-�Vm���K�x�[��ַ5�C�o��u�	n�����7�|SL|�Yo��.��~�w�$.u6ێ����K%F�⺕0��r�M��`��VY<Sk�Z
6D��u�._��Lۀ�ME��7�b��4�o����{�?Y�J���WM�N������^.i^�Y7Y2¾v�Zuaq�#ZX�Z2A��Z�����o��ۙ�"��Jn��a��bJ��i�W��˫�JS�X���,��<�`�aY�Rcso��x�t������ ���hw�,S�lӊ�$����fI��=��*�C�ب�h�&]�a�-LŻ>\+���N�o8i�5�ȁV�I%I�����"FS���ܳ������Rl;��[�R�{���m��+�0��C��f���)S>��gd�Tl�V��l�J+�_W>O���gY���βYٹsn5� .�����@���xJ4�� �vؓ^�D���*ⓔQ������dY�� ����#�Eĺ�T��Ņ~8ren��[��H�M���Z\׷]�rd��]d�<�)!����0�,v\��`Z��������5b%;v/��J��ȝ~o;�� ,3�
�l4ԫ5|��h\����7�ʶ/��r<I_dc>��/.-�����p�ǳ]�<�z�Y�u��������������7ĭ���~��Q��.�15��U9�0z�w7.^��K/9�v�؁��eب]��[��R�>��93��&G�t:f��+���;�{A�;q���Bk8��>�h��G����~_���<�[45�T�����6̀�j,��8��6>�-K�0Y����i~aae��=����~��/ի�F��Y�2\^Dy1��ģ��4_b��IʠLo��O�s$��ްa�{����~�����L.�'���¾�"&<���`a{�t.�$T��0�W/owol�n�T���p9�|O� ��j@��H���)���G���
c��-ee �xt�4ͱ�|jr�![���(�-�,�| ^!+<#���?�G��BN��������١Ga���P�E��d�Z0�-�j�N��>.&#�dL�>�4ԁwJi��k�O/·@,��\V8�s��勣�զX�5�u*0��n�6�C8�x��i�Nb�5��E�uC�_���+��%����>4}
�����X����e�^&O"��#�iO�N�`y�W��Zs2G �HE(R8]��Z���z{i-�����_l��x��w/]���c;z�(^�x0t+#�$L~ ��hf�n������a��W���Ry�;4�*�w��/�~;:����j�[/}3#�(����N#s)/��7�E��Y<j�#��I�"��[�ݜ��_�u|q0
�W3u�p��C&�����K�;��k\c����<�����2<� �⌦�RǢz����,�Tec�6�y�ӕD�3@���2�{)9��b�͖D���Z�>����R�4:�y��$q�TLUS:��-珌(�M��ksk�b3{�;C���*1�������(��v�]|�3 ~q�,����Sa&Za�(�W�΢^vj�T���z��g��1�{�/�Bc�wr5#Zɗ�bj���fz�9J�Pi�;��ȓس���E½�
�N"�H�����/�?��<ә!E3��nWn(*'��N��R�0DO�}ْ����:�VǳtO;�0	EȊ�+âb,sm��/�>i�#C�ڔ��!b	3e�r戋Y�!���m�X��G��+�b�k���Y\\Dd�~dhT@��Ջ��Ǳ�uggOye*�lΛii��I/�,�T�(׈�M�}�����A�(-��G���0����қTBq�����uL�t����:̲G>�|HJ�mW������\��p.>�:�)�,u:��ׯ�ٸ޸I�&�Ql��E��Y�//�`alߺK�ϤɸR ��;=Ɇ;�Q>�E�L�Lj޸�u���Z}������5{��h��D�'wc��������~�b}��K��1Z�gZ�=sx�T�P�f��m�{�z��7���,��QF�P�v�e��(ç�R3SC��9K��{Q���uRx/�%��L���ɶG�Ybp�2��e�(��d��gfgDF(��f�':���?ˤ@+����y�=���<����j�J��r�8�#ؼ,{�hy�ԦL�w��$!ׯ0ݾ�����K�y��w����T��Γ��8�o2F��v�?���Zfb�1m΁W�FZX�8��]�&&�S*�<�As�eGN�\f�e�u�^9xՠ��gv���L�J�>�KC�z�A�Ͳ�c�4�g~��1�qY�TբaɅ�^o�����%�U��Yia��iTF��b�բ�5X�QE;�#�π�:l88�5<��Ҳ���u�Wx>rx��&����9?&�u~9�)���bȅqEq��q
���S��ŋ'�e�4Q�-5����2zZ+Sq-�(��f��9>dB>�Da^�Jf���*dh*W��xr��p
#x�z��\�ƭh�@�Wؘ��T�(�֪�f�1���]9�9a����M[s�� ��zVog{wgn}ݩ�At���+����?-�
̠��+�VV����/�|ks[ľΞ������֖WW<|�
��*�A�ƵO�a٠��6k�:)%Q5���`���q�ȑ7���7��MW�&��~��#M��Z�My#�gM�|�e��^�'��F����(�Y�zxe����J�62Z�D���)�8���p]L���c����J	{nyVA�%��ԫT�·$ߺy�5W��`gɢB�4ES$c)�玎c��-�m�#��p[�L7j���}
�/1MP�;�j�c�}H
A�np��i�����0Ѥ���>�M�˕��Ir�� H�7+���h�3_
\jg���/7����A�tĴ����o68{w�՞[�a`w���^����L�oa8k�nN�`�y﷛$ULl:�S�E���
��K9e������&*���1:9�{A[���2�".�7�5��A2�����]�����=���\�R�S ��1���<�Ŋ�m�9ǎY-D+'��m{{�����z���W�^q�0���	ez�/L|J<��X�V�Յ��u�SА�C)?\�}+?�Ke��(����GÑ��:�o���~�i�����ţ���	��*�ㅙ����J�>��D�آ".�y���BW>
k���ǟ������\˖�4��) "I�� ;Ұ>y �d��qxN8��5�Y�Ƿ[K�+�8����4���O�8�]xc�6aF��8M���]��6$�]�^3@�x�닦Ή��o1����s��(�%��˽ �	�H�����hx�5L���ˬ��������^�sp�;>��@�Xo���~�K �XivR��	�N��0�2ܟ+l+��ȍ�,��{Կ�G-�K:'ք_& #���b�"j�c+����&q�R٥ԋk穒(&�3.Yʘ����(����g�$��p����;ר�A�i�dd��Ж��h�M�J�Xƹ��R���L2�Ǽi%��l[��ȍ�|R�t�!�[�>�[�(�v�Q2��l�"���CS{'rrByBt�〶S0'�9�8G<�vv7n�x`�숴��@\X���`<"�E�p�o0�DG� �jo��� ��	4�<2�>�v����B��}G�� P�e���YE��U.��$2q��\&em3U�i�<�5@y��ֵ��3|n�д𥾟Y+�"��!�(r& ��S�v�*VdhKX�"��W�)�=��)�@�>(z\f�O����	ztf��xפ�[��3�yLH��	���	 ��N�B�i��I�$.'VH�S�9b3�����~�/M��mev>Rf�q͘���H!*���Z�w���v Y8`�������'VV��%�xqy5O��ht��C�x��׮\���X8u���B���M|�Q��_�=�v�m���nD2m�Ǻ<�蓟���'�}i������Ϯ�nm���{��]����/,m���z���T���G�\���;N��l_x�V8�u���C�p\�v5
a+����`���L\�Y�a�;y�Nd�����i� �l��;tg|��u�,*α�c,&��e
�w�*�Ғ��L��n�G��B??��:������U0C&�L�Q�n������^��ٙx8�ne����P��iyyykk�e^N�*�?���DA�+�f��БȞ��P�Z��~`m<��t)p��A(d$�4�M��o�v>)��4u}?��f�����6pO���KF3	v�4���9O&�h↑(S-�j�P�C-�n�k6�o�BclVj8�`���_k5o<��_�z��Դ]l�>��Yq;yh�6\y����ue����[�3��I;4�Uj�~?40R(d������ӪW#S��B���)v�8$KN��A��� ^V<N����5d�تW֗W�����{�v:,u(�$Ê����8M���V+~�uJ���cm0��Z�Rca�%<|c�I�Ke�X��ȨVvvv�J���nw�'�?c�O�Y� � �?2'�Zk/+MY�@�j��Z���'�EA�\'�`�f�p�;S�u�rsi�񌰁J��-�S7+�#2 K�`M�p���9^�*CL���� ^��>1$іy�ڀ���}7���j N�A8ߪ[���飭N3�7MBCTuj��U�L���$V�t�H���h4�ôV��`~`�2K��qw&���:�A�J �Zi�$c�wnЏ�O�D:� ��8�Uw�{���k�?@F�#
`��h��j_�E�1�`�/t*���D�C/w
�?I-ȱ�~��ְ�?�O��R-����C�~f���D�&����
�h���M�/��E�8�md��%�'if��2o��h�-8FP�C���ܾO^'��Y�"�@��^�δ�-�⻁o�aè�A��V��n��LEI��>��(,M�S�ܱt{�z˫:i��$�o�D~j8�VT����L�� Șt�&�T4�G�_p}}]x&���ʊ̸�!��|����Ｌb�0Z��2YnF<GI�3v�L�.knN�'���4�r�#~���L�Ih�{ʇ��wk�֔�
�3������/y:�V��mEte��>����y2:�\vת��2!P��˗G@HT�|���:
I�W
�(�'	�љ�'�����3c�]@J!�#�t���9���)��?�8�Z�wJ'J��d6�/3�lO��N��s�æ�$����xJ�'���4��dX�Τ�X��?E���i�)A�i	����L�"+����8uw��6o!�\_[{��ǎ^�t��k׮�^���Ro6�\;��6臷�U����kw��9����ϟ�r���ͽť�3g�6�q��tqc{��i�;�k׮\�t	��+"Hg[� ���e�N616w�UYO�q����?N:>�_���
۾5���F+�➍����Z*�2K�q	�?� M�/T��o-3�F������H��M�,�)'�3�~���&\Q�n��\�o0-�cAA5�Rify���+�;:#Ǟ��s4����I}-�ޯXQ�����e~����-:��lh�Ԟ�#^.ɋA�Z��?��'�|ҵe���'kM���K�8>r��;��\Γ��#�f����_ZZ�5x����N�>�Slo�bў9sfaa�{uu��p��`<�'|�{��U�x�8�>�y��j�պ����'���xY�q�Nt��ɬp�������W�T�"��Kz����:�����76D�HHeu8GՊІҲ}VV3�N��=�g��>M�i���t��=v:. �%�sf��&��i�@�=z�nww���.$8a'a��ǅGg��2�әJx�D�}t97A��M�+H�v��0�U·���f��4�ƴ��1�����>B��<^\\�:'p��{��c��^����ܺ��r��H�Q՜ۖ'�~���Jk�r����$y4�m�Vo��������E����` ���<'�BխX���`��H2�IQ��j����C���w<��$$B���Qh��\ӏ�ync�r[�¼��{{R�v�+�M7X=�̵:c��[�]3�1�W	Z����J���v���@Tg�T���mmm�g:��ec����2����1S=M��d�g!�?�t�r��ǐ"|����9����]%��pw�L�כbz��]8��\:��𬱛E�=�S�e�=�I�<ʢ4�澗��Q�S�9�Y����H�)��\)[%�2��w��0�&�cc��8�M��5�{L�>�tr�b�s�&���&�(e��B.�.��v`�)m!��ܡ�=m�T�HYS-]9*ґ�eEN��3�ՌuY���8@==�Oi�Ud�l��h5CA- k	L���S�	f\�^���L7���+��&�fߙ<��":5Ue�a�y��Qn�����3����:U�X�)������)@*G�)R�SM᳓^��M���3�/��t�ߦr�%�U�]��j�Go��|"^،܂!r<aӔ��5	�����é��x��(s�_1���!�ct�-.�p[��ml޸���?������n6._���;o��¹G[^]iV��4�u�7v�v�0�ӏ=��;���W_����;����s���no�?�I�����q�z�O������f����Ν4�l���&�i�K�f���mͶ��3��J�v���P��Y�d�x6߭�2Y$w���IUr���)�Y���e�@~�mPtG3	-�m�N#ϕ6Q��f��ng�Pf���_�L��C8����+��f�jc� ����R1S0�W�Je�c-�߳Y���׻�m8Ӊ^~�̩���<7�4�N�� �Xd��(L?�����/�wO=��4��E��2�QL�MT�ޠ�%q��vl`�m
Q"��Y�|U�zE��
0~�u��;;;�����$�-9B8aF`�"ˁ�$Q"�Wj��-3%�� ��Y�, �3j����8��c����.N��������/�3�#�A�ƙ�J�[f��9U\EMc�D�a�|>W�����K�D�'�=nh�cU��ʅ%�Ճ)��6N���.�O-���~��)�aa�&���Oy�Py�k����dx����R���3��2�����,c�<BG�PnGssK솢�*��@;0�Fw�Ú���[vǩ�Ii~�$:��5�p�=R�!��F�p1�F����Q����_��׾��hiq.�ǣ})�! ����^F��s�����ԫ��ᙩ<R����ص��v�^k�{2�
ǜv�� E��툵FDX5$��s�'�B�ՂʡCk����=��+++x2����R=s�F�9�0_}䑽흫W��X�FY�=U5�I��;?om��{�͛�W/_���?�ܼy�?Lk�|g{cqi�#�s�.�ɲ*D���1�!:x�'L�LZH�I��lq�1����ӊ�}�c���
���pA�Ĳ�S)r�>��*�69l�h���4L�p�ϭ�S�LV���"q�QRV�,�a;��,S���:���!++Ea�;�von�ˌ����8�:�<7��7��2�c�m�rӉ�I@��7��<x�>W�u�����w�M8�zK��0Ӈ]Β�E{��&�GD�>��|{�"��T�Z1%�1��UpU6�,ш(�MC�r���*O��53,��{�ʲlJY�6�F*G"rY�n澬Ҝ;m�b�l�{��0����� �L�t�J(�S�	�N��D̡IwT�H���-�b
�H{S%%�J��S.�i"�\���^� 8a:�
���b3"�����P��hWmns?�N����SV�uk�N����%�C��WI��ygg֮Q�Ê�敪��w_��w���~�~��Tͭ��o��΍K���WϜ{|�Z��^<�b�wiq����Nnk	�E�:�wӴ�D�"�oy��h����5mf��J͑�J�6uː��~��ۅ�8��f���vvn��ҋ��]w8��w�����{�j�=����L��~�T��7�&*��_�F_٢�����g�$5E��DE�V�sa�n�yiW3��`��?��Q�B��R�AN�jn�L�����X�S���Be?d���g�2����m}xO���
Xw��LgF��:�F�� 2��]�6T33"�qp��I��?\��7i��m��a�#c�e�Rj���{�\���X���v�X��y��eIf��+벭���ŵB�nI��h{�����u:J3�`���fؓ����2��8L��+�3����1sᖳ<s��?��s_~��W�5�^�J�&�����v������<V�<��>�T<��(�\��&���:K�����7SI��q��"'G����q���>� �ǘɄ-$P0�HfN��߸qC�
�g��3k��O��АZ%}mzj\!�Lp:�|Fٵ��f�#�T� _�ˆ(-yu����ld;v�СClvŽ�:����Q�W�A^*g���4K[L!36���$�|�Dy��F�G�~�'rp�k{{����W~�גxT����N�|��Y��#�ۍ��9��~������3�(~�2�p�<� �Ngaww��ի�\��F��K�\�܀P�`;��i"R.���D�Ï�����?��c�Vxo��Ƌ/�x��%�cD�[۷�S�N\?�_t��˗.햕g���Օ���b�Ҙ�,�/�|��׿{����V���<���|��l�lu���j�'��f���^B	�5oZ�1T]Y*d�Y�AH�Ֆ8$Q��'F]���i���4�:3��|r�I�΀�������/E'*�� ���#6Us�;E\d�D�j�YX�#�Ѿ���a�R7+��H�ٳ*k�)"��b��Q��=@Ң�̖��ǹF.���������g˰�ƴ��9�Qn��*>�ff���s;a�n�!�����v��(�V���R�إ���tX��e�
��Z�¥�oZ�*X��:�Z� �(��ZBaį_/w@)\�8C���hZ�t��+��!���,�TFkeѼ�����ɔ�*B1�+zt���������G�D�j:�̣��Δ��3�d�C�>Q浼H���:��E�K4�W� 
()��U	P�SY�H�����u�q�g�0�C�~����/-=��
ana��l�����>ck����?Uk��n��N���t{{�Μ�;?�3�~�����	���-�3�O{�Әk]�����gZ[;�z�j���Q<���|ggo��������>�����������wq�Y����ҷLaq�����r��W�W�G���l;����)��'�2��b�sU��̠���~&0*/l��V���D57�&�><�7k&������ض��8M�|��X*����s�$�Q4�j��8���}�c����u郫[[[,�r��?�`���@����h*�iK�:�}3��|���&��z�.I �h�omn��/E�t�;�`Q���M|4�d�#D����5Jr3Œ��N��h[�c��(q�5#~���$����D+�^k6��nw7
��$�W�����V��#������*N�ͬ4w�$�#��W�Ǆ��Zs�}��O= $���}D���M�s1�<����"�$^������|�J�S�K�1��KKK�#>LO<�+W� �g��,���0���a=�&OJ&�bQ��$ʄ�[�&?�nh�Q+-3Ɉr�b )ݔ�m��YH��3��u9�V�0ޝ0-]��_QƩ�8q�����í[;���D�ՈM��\P�gsM}`\�e�O��06MK���!c����j�m��J4ƣ6��Y���xwg<�\x�����ebU��y���=��W���?��?9��3��[Z��J^X�����
l���t��K����;	2���$��1�&�%1��Gq��̳�9r�Y�^o[���3'��(
����8lTk��Ci$
�J5��E�������Kqj���Q������̃����/{���V�C��|~f�E~Y���4sHtG�4�I8"o��s�Hb:��I��ɀ��$��`�:�B�6c��`��8�>�$�X8y�c�q&���{�ؠ+I��U�"M"l��zn�}��#����iq �@#W*98>�2���G�nlx����?��!I�b� QL��L�I�S�T]wE�/m��T}?�N�$�D�;�t�S�L��#�2*�%m�,S��~]iW�@������#jcu�ͨ�����P[zڈ�l&��:�@;��>@X�����#�c$�� h�ge�k�����O��*�tO��8�C��HSQ��-��B$����+G������xS3#S�YFw�TƄ��sOj"����d=��24�%�W/�ߝ���^����.��ݵ5H��j�+lֿ����eB�sHq�G��/C�j�v��`"�[�p�o0
��3������a�'V�	4�lo O@��oa�}��Ϭ����o�~���gϝ{�����ե�>6v84��Ȳ[��*�:���\�i9~�xn��Π��ks�x���/$�������B%����<��A��[�l�ܺg���>��*+$\���j�� ��u����i�k����<)��{F�wS���)����^�t��M�Fbn��	�����̬�;ڂ�O1e�I�p1�|�36���:%���&�0�{�>���onm!�=~�8�. B� #7�`0d�~�Wև̸�J��3�����r�}���Xx'��~WY3S&�l�Ͱ����|!�.v�9�}��o�r���F��lց�;�ݮh�̵��q���@�Pf�:`�JS�1�P���7��8�������͛�G�~f��������ի�Q�=8�l���y<|�K��\�eo��׬�H����1�aT�j���/4�s�Z%����ǟ~z��l�QG���:Z���VV��;�T�!�U�x�W�&�yi�doF�\���=�裿�����#������/�_��H��O��L�.�8������p�B$?E�K��n����_���I�G���d'*ٔ3h�ՙ��̘���IegD@�*���T�Q�M�%�_Mx&cՓ��X�ݽ���������/�Aq��Cr�͛7N�:m�Gu�����hd��v��h�C���Q����������s�-��D<��$���G��x����3g��7����ޝ_� X96��b����G�:t����������W��O<y��������^���a�ܹ�>���7�_� ����1�s��^O�A
�1Y�$�s�w�2>s�ʵ���"� ^��?�yΩN�~�`�(DT�Vwǣ�͛�ׯƣa�Y?q�H��Q��>��ǟ�����+.�5��U<��cG?B>� B�f��UI�JR)3*����k|�H���[2�{��{�Ĳ�e2-����-�v-��p�}��a�ѱv��P��*|�a������n��(��N6<iؔBP��=Ѥ�t��m�@�\����eO������@D®��ĠL'�y2*$+D#����f[egdU�����///�{;x)�_��q}}m���]�8;������cX�µ�5��23-����)AY���y+���es�<4�����BE�h|�E��\�tN�9��U{�\�Wn��q6�6A�Z����t�:l[�3�G!�5xʂ�|�2�芈s�x��M~JHS� �*�F̣ @/�i�[��w�ËQ�rͰ\ښ�bRjfa�lG�����~T�S.^�!�72�K1#�W��-_a��g��a�,���\�v�?^ZZ��&�!�c�,+��<I�F����"�K�R���{Y��� ��>��c��/=��kgN>�Ѓ�c�N���ي��>xp�8�Yt��w�|�ukGO��7�v�X˪՛�}����y}[�I*j������|���ϟ��7�y�B�lک0���2��u�"�����AOPnRܻ��M�9FR3�m�O�n���g��Lp!��̈v8��kY��t_���V�"���4�/��k�v3�Ԇض=��px�f�H`2�cұ$�Cn��z!��~�ۯ����H���6-�Nʡb�˝<�� �_���f�{�~�r1�l�gz5�9堚�Ia0	h���o��Ea����ި�s���N�W��_�����'� �T�����n��]wΤw��S��Ep/��*8;5�/�q׮]��
�UrɤU`J�*v��(hTh��$�Y�����ے5�j�F0���רW�Qx��c�>���f2�Cڞ��������#͆�Z��|���߁Y�t:��qU�T����{���Nj��+ģI:cn�����x����a�!L�{��w/^�$�vm}	�3.`�ڵk7���������{���l .���~���v����ńT6�\ *ﻻkA�V˃Pu�����3Z�Wr(t��l�w(d��v���W��ɉ�G�����T���W.������RL��j�����'?�Ƀ9r��iqF|�<�?����M637�;�~@A��B��y��_���6�q=;���pԨ7+��sk0܏�����ť�j���k��ny���ھ�������ij��vw{�_[[:v��8޺�y��e\�c{y�Q{.Ax�^��ʲ�7s��6�a��\Ey����W��_?w�a,�˗/�E�ƱN�I��UX�{��ဓ�q1�����1��� n��,�,�;d��\D�f�n���7�Gi��9F����@U�I"31��c+NM"M�
2��4������穡���&3�>T��.�C�_)��%�b�pk��fv�aw?�F���zi�8^aW	cS�Q��N����N�`��hK�qBdrR"��(\+��v���/mB��N����^ھ�]Y�{��*�oI	$�I��	{dcs
�Sũ9&4Wn�:Q�6�ra�)���o-�(����f�T%���t�Tv�V2�ԩ������H;*x2VV$�{�XA�6ю`�xl*���NF2/���J����I�(�pK�3��)[�$�N#'�Gq;.����=*��Lq�#,�����[���$��˥<,H���9BXO�'"b�,5�Д�0	���Tf8(ޛ��MA�gڨS�l�u-�u��B3�|�P�����qj�V��Yܛi�(˾�����H�伮�h�Z��zoow�֦���*�Z���Agw/�0
Nf
n'�Q��|����`kAu�;��_~����N��G�7�5�Wl'��7N�:?3���X��/bDQ�F�nŗ�H�?���8���x��awGY͌�y���~�?�DQ�0�M���!�������7bo����ٰ���՛\������W���X��87��I��p^kv��L���;]�&�!���Lu�i�6�rR�2z� ���i;���|�&���܃8�ĨV*�j%��rBdY~(��4�)#��bQ.��`�V�LE�C��@H��ʪ�����2��&Q������7���`��<�w{W.�:���+��B���-��s��#jW�Mv���� 2���M�KU$jO�p�%c` ��a_$���DuX�A?� aڕ�0�Y�ا?���j;����C���k�g6���`�Qs�0��]uݴ�?����ׁ��Ү�Zqb������Յ��č�`^8��g�凼��<��+����1#tm�7C���(pBS�f~Ξ=�P$�q�ӧOS� ��^{뭷:��?��C��p�s�Z�1��C�o����z�*�����K_��A�M���t�m�i�����n��Uޛ$D�t�~):�j�Viڵ']��ݘ�Sm^�t�Q�����C�1*p����ss�����n����/����|fii	0 �����@�ԩS���g����r��Μ~��dW��/=i>�4�?�d|�O�Ӭ�I��[oy��f��p�چߏ�1���#G�xⱕ�U��>�q��g#2	k��~�v����EY����>t�����￷��US�2����aG��:G�/�Py0����}�O�x�\�����g����$1]k�ۍ���¹ӧ���"���f�qG���bg�רׂJPC��d�}���h��V<�5�p�D�?�vGT���Q��\��,4 �#�:�Y��2�ͱ*X��es����NR�Qޢβ�f���'5J��RI/fr�f��	XEht8�')@���i�Z2��I�^��zF ́o�t(+L�iH�#ͱO��������+����-!�L��ovl/�Ճ�h0�'����`p(��o�E��"�����N�gg��9�-��B�ǅ�dK8nKt�+��a�Q@&�Ņ�/&�Á4��Q��%�d�a:�O��Q����1�-P���q-�������a�Yqd�c������ډ=w&Y4f����5����eiE#U��e'��ж,�Pn�ц~:l�epi0Ę���IZӜ(�/�E��q-ώ���1�L?c�+|��'`��ؑ=��P����L��K����F�&&������1�2Y񀽃�����B\��˗�E�P$Á�*DԘ>z�(N��������_ǁ5Ƿ�(�@�p��$� �Nt����Ph�?��p/2mwa���:C%���{��¿2K`�Gʡ"�!��Dz�.���5>mY�%d�`�	P����G������QQ��@�ZR/H������Y���$���1<d��)��@U�T�N����0	^��V����/{�f0�E��������ClC�L�o�-T�V����s���<Z]\D�9ڸy���"�J}m���⺤{���7��ݥ�ΰ�ը6^�c����x0��Ul��q�Y��Z�^_�1���k����J]�J�M�N���R�Yn�e���]`Q�nܬ���#;^,���D���fAf���ꍎVd��5�eF�u�!�M��$̐��fbW��T"�[cp�Ԉ4��<������ ��J�Q{��ĉ/t�Icc�� 3��]��5��\���k�p4m�)�a���ar
	�B8��	qIB��Ҵ�[�@�Zz���F��Ε,r�wf�K=Q�~�����:��q��&��4�ԑ\���ԦMnua	�G�jZ$�Պ��l�
��{������T��P=s���vv�vejP>�ܺ�����G�(.�xs�^�v�e�Һp�r���>��\��/
i�j�Z�{�\_-���h�ì]�j�Nw�ԩ�����'<w��������ys����W����27?���8��	�S֜���Uq�`���u"Y�Nx��Zŋ;tH�"��L𛦍�&t)��i�� X���?v�p�Q�ޛ�͢h��pl� ����y����s��Ix"��d:�Z��_n6�gϜ�,/��D�f�c���$�Ç�+���'^z�K�.�&3H�E�N��aAe�V�ŻU|t��O*j2��r�ic*���
T|�5Fkϣi_�	����_��������Y�Ґ��R��w����x�)��~�'��hƒf���`�W��X�P�(�-_.zY�%�	��DVa�$�l��R��2��jE�Nn|�Xn��ĩ���v�رg�ӕJ��?�p�ʍ��0�#��8J}qCNg�q��i���7��(��(d�U��k^�8���u�S��ׯl���­��ܸ�}���=����hI:^Xlϛ�U4i�����{�&K��Z0}�嫺��n�A7� A��IQO�PL���}�Ǚ�0�E�?I��<#�(Z� ��k4�޻�r]�����Y��NT7 P�o�"�y�V��'��{�m֖�B����*+�ACr7<����f�f�Y����.U�L�l�%��������	��X���F�řoY;ggv��_8�or�KÞc����o$Nr�[$(�#�l!���=��p����ڍ5���9C�8�٨�z���vś��dCfx��$5�	[�sO��aw��`{;n��I6L��E!�!SZ-����SNw1� ��sĖ2
�Q?|hn�������5Qo4�����$����[���tT~�=�a0��mg�lT+�f32�L����t!6�f}ԥ J �`�����%Q4ʣ�I�!{�V<���O#�ެiAY�P���RƱl]�c���V����~���f�kO���b��Z��q0}�0
bۡX��� �pZ�/f����8��� i`�����ĉ�'O^�t�ڵk�& ̹s�H�
	[�����ѣGq$P�|����ׯ����-��b �J$���ׇ��U���7$?X��p�fffΞ=#=4�͏>��-h1$|��믟:ujaa�g?��ÇO�>�G��>�~T��#<����rq5|օ�X�9�ǘ1��;wb08 �Y��^�i�u Ҡ�y`<c���X]@A����Y+��1o,��E^z�%<~�eɨK�W6���*#Ư�O��..�,����e�1*�J���L�w���S�A��� `��t�M��0�4�vXLh���m[�����m �x��R��BȬ��¶�]^x� (E��s��,���e1>%�B:�ޡC|Xu[k��k�FVo��~�F��Rζ���Xi��MOOa���֮]�Zccw����t��5�������S5�f#�%R�tÝn�����K��~��UQ�N�<ڶ:���L�?�"�j�����W�j��[8�LR'kVb�Ib�`��X,z�\�l���?�]�Y��Bُy�4�L��&�QI�B��D��X��7����4�����fqbb��� ~��=$n��V����R�F��9~��?�/��k�����8�s{"=k��P��i��Bqm3��'*˘�V! �����$�`K���͗�z����;w��t�!W�^�-�Ee�����8d����3gO��G�����o���_��_��d�è��8�p �eab1ؒ�T��9����?������~��m8������ǰZ,Sj���O�����I��:W�^���;.�67��Yy���������/2J<����H�)�g4�d"�&<+[y�K@�'�WA�V�{���S�jw��!a��4���3jXGwKS�zmHx�m�o�|H�����:z\�aӚ�JV/~]���N�*@��������z;=�f��Puu�a�^�ܮ��Q�ـB�CgA#��3F�^:O��!5<K���������_e|��R'ŐI\څ�!���]���u��Cha�Tt=�L�$�)%�f�y��=���* �ZbTݕ�kW#a`�ۣ�ᰡ��#H�T8#O���#�CH+Hy.�%1���fg�xL�D��ҕd���O��m�*����S@�X4+3�rU!�f)�z����_=�pnb,�m-=YZ��>�����+��a94�����*���[�ꊇ Z��ڭNo�tl5�X	�Kk����Ԛ�@^���"wr��f�U�kBa�$�`ss}s�cc����&9��2WE Eq�k�<VXQf���z�.L���)��t�m,,�8���ZKx/��5��!�-�0�̳K��$�߰M#�%7=!i[lK�����n�j,�pk���;V�Pm�?��A��\��[��X|0��f+ӄl�7��)#1�F��D��u`'KC�*�4�6"5~4��6~m]��9t�7:���o���#��T�q�]t�2Q^u���5�Rx�"�Gz�0	�97]�@�:��/�]s ��5a�*�nX�W�^����r�
4 ��9<�� `�+�ИAe ���Yp8��o`��.����qLiy13���\�/��|@�%x
�0o߾|ŀ��h�F�-8�XҰ����e���\�G�GT��뼶�[` w�������x|�O�+��n~��1��4;H|��Y����g�ַ�H�s�U�h?Q?�2S)0H��k_����c�����ğ��o|��_�tAjC�c�y�w���xL;���� \��[o�h69�.#$a �
�N�ԙ�A�A����,A����������zjj@��<�J,�JqC�.J
e�ܜeQ�~s�Z���6�&�g]�k�k� B�F�@L|�LO��`�?|x�����s�~�۷wo{r�ڥK]�p�=��4k�c�<4� k�ډS/`�?��9�	T�jt�+���Q5n�v�V���Sۚ�|�%�=�pV�ab�0;�4��Ma�U�ط/��ٞm_��1��j�؊��'���3�`��㭫:�ua h��5���(���1�4�[��=+�q��~@��I3��-P�u+�s�ݻ3�cn��t^.��[lk��-G�UF�b�j�P=-3��eU	NĒ��@��2�4�b�`a��$��G������f�Yn�~���>�t��=@������a��.'}��{����ԅ�]��%t�L�x��ļ
�كA�^o�9���Z;w�����j^�Ɛ�8���,�����9�-X�,.=�˿h`�nnn͍��g;}M��.�����7�3�w����Y=v��l.i������k#��tlS��T����̜j�wR}ւ�r:�BF;D&�x
���.�V�6F֪O�+A��?͔�<��򨫘j���=A�eS㶑��~�biX2�7Y�C�-Q茶���ό���MLO٪宦�ħ�pW2�oa��	E/��P��Oո-Ö��Ȑi�wпP���o߾����,?Hxx+I��3'_<�c~�,������m�J��(��y}}F)7�L��W�!N���.��$�B�Ʋ�
2���#ϟ�
����$Y���,4ۻ�=;��Q�/a��E�LK�
�v�����������釯��Yׯ^\\�aYX�V)~$��`4� ʾ�n��'�S�Y�@���4
?�F?�����|�fR5>q�Mk���be@�Î�6�<���*�
��Cf�I	���eV�i��d[��L��F[9��ԓ��L�z|���V�0�6{In�ON$��;"��V�^|�/ݚ�II]n+��ϒ ��� ��"��T=ׂdT��©�&!-lR�sS�2ۃ*8Wm����ؙì�QeKi�(������)!ZI#S�Y�X�SpU�;׊�Y���]�h��jH��J����!��J��V��<�M{��tZ��\�?P�ÃYC�m)]�Y�跃�M��B��{��ě7ob�`��Ԗ����C"�Wr� ܹs��љ^��Mh/\���ώ���]0�3g���F�1���+���|��G_<�l��i��a�׋/��+�������4�/_��?���.\����;�����4���W� @,N���������E��qS�.�e�x���GrX���$��Q�ΌA<��㦘I��0WxX�]�0�� ��B���1��<���W̃ϸ����Sۮ� |����X�L�(�����9�1%BnE� >d���G�.���s1<i\>6��ƽ�wp;%�"{��!�ΑV�A݇�76�:��ɫ�����/�<�hbw�y0(���֞l�L�2MS���0�,�	b�0��76ffw�]�]�vun^�dCE�`A~�?����aA�w���TML����t�F�V�9ڑ�4�jE�g��TZ PUc�����:o�,]�M�=L,�<_2m�J��Y�5��W-�t#$s>I@��5�~��]��8
_��XN���� SSx��+�$�*�#�k��e%��^��ƺQ�<5��A�ᲧO��=||���MEC����V״mEG�6O[���C���2����̓��$�a/]H�nܗ.��}�չ����b(273��p�v�9�w��۷nܼz���0Da�������?��^��N�`6�e/��`�(6��ʪmA�{>�pcmX�,�,��鹉��Hj~��E!Y[�J������N������|�W����OQo�(R]��������VXE۪e��4L���75?,2�^�$u��;X�#��r�����ip�8�a���)�(iп�+@�+Tu�y��G��uׇm��k�D[k|]�>tu��Yw����d�!��Ӑc��U5���~Sa-�U)�<eJT{P��R]]}=���R�z�:�:�S6/X�5�9��2]���?�/^ܸ�l����ZP���  :���%AA�����Q��wO���	Q w
�Q�V<mA�1�~���q���3U����%���ע��<���������X��R/L��H���ύ����Ŀ�����NN|�;�3���wh���������s_9���~����w���oߊ�pj|�ccu�ӭ��2�����6��f�c�waHg9�;�t�(�3\�Q� �f�t����U���NQ������~��rӍSHa��"+�����b����r����XQbH~IOr+q_���f��6� 6��&@6�Y��'�B-��L]�[�C�C!b4IR�)J��uBCf�σC41��S�F�T䶶��1t�U�Lg dЎ��H�$��Ӆe"a�nHF�ͰN΍�9��6�<�5�:D��Aլ-t�L��4V(�u�����82��v~T)�hW�x� ї�d9!h{�t�:��%;#Qǀ�I�|�$ZK��V2�]�vI��;0����Ò�޻�G ��S���2�z�j�P�	F�2Υ���� f�\���8�޽{��ѣG�)+��ɓ�+�'�`z7�˹s�10l\AW@qn�h�@��10�z�a�[��������瓸�;＃s9!+++�F�zL,ln����k�Ξ=��%bN&�1��``��w��]�������ZXX���\���
]�|eԬ�#q IF8��Ǘ@���`0�T$GbQS���̳̇�]�,HMm��:x�^�����P�q���C��1ጌ�Y�B���X{�����������W�]���i���y�-Է��;u�����;kI�{scc��w`I]�����d�asb|ffNvh*��x�O�\�W�f���z?����]��W�0rU%����'�/K���V�(��ی`�b&jnK0{��ȶ�����Ak�ju�0bo�R�����[���,�%0<IOOG���,6	�֨^m�|N�^U��0�0�ESd�ǿ�e�.��}�~���;v�0.�w�a ��`a!�$61p��z0W�^�L�9N1</ �9@ｻ:�= ʎ1�[�v��T5&�,k�P�_����!�OcK<ʑt���ɣ,��L�X��<|���4���a�=~����M_Y��;��?p��ę3�F�Ⴥť��F�97}���z�na/w6(̛��V���:�L��j,,ޙ�������߳k������^������8%%�� V
S�a���=z�4��)O�m5��VgLEuL�2�[���S�ԍ%9�c#̖�$�*nbr_V���iz�&0u�D��G�LLLa�cb���4�A]��s���Q�#��u��Ym4ϐ�η��P�Uy55'�SQa���MWC%:��{��a�l��*�n-t��x?�4DQ�n�Ҁ�SlP�av1��k0���ge,�Ku�� �C
������v����&U%��,WS�����Տ쁻�����NRe��n'�}����=�k�Π6�Ձ!'ToE�a6}o�<�,���y&��*ĈYpP���Bw�P��;���4��q�	��8���0s���0��B�>�R�M!=��纴�CZ�/1�g!Sr�l,/�,�^���:tl��|�������d����X`X[�^T�Aq0����L�� �zP�e&}��H��K��@j{|�c��&}�T�����I�C�@�rSY�
T��[�K��n؎�v�;H��Ȝ�i���7ղ��8Gb��pٖ��2����1n�[�U��c�z{�7TR���p��O���^R�9y��;\���Ryn3�O��(Q��̚2�|_V�1n[��Vw쮴-����:>%���r�F�MW8m��~�m&�P�c5?�C���tn�-�f3W�c;��Q�u�pS��݋��b���P��U׬6�5���2�����:�d�]��y�=�!5Z9�Չ���H�X<L��t#����ŀu�M�0!�s���߰�����w�Իo|�4�9`�þN ���Æ����e>q��lD�JHXz���' B��.��א]�1ƦΜ9Y���-�rU�s����q<�~���4�Pi֡R�0$�0l:)�{���Y��p֡wݼy�ez! &`<w�ޅ^�ɡD}����&� ����1qAsE�8��q��Q���k�w�e�<���Ӏ�x�w�9��rC/l�#��*�}�1.���'��xo�.	l�v�,�s%ب_�r�p�c'άl����[ᑓ'�4ZYX�՚{v�3������޽���6j��n6u��O../CjP��_��л��^<y�y��MY����� ���y5+���j�m�E�+�$��<Z�?[����t#c�t0'���*� ��ŋ�?,`�"�����fj�f��V��hL�O� A8=�M��.�I���wG�z6����Ϣm�C���ع{g�7���t�6.6���+P]���@�i�Ƨ;U���
����Ug�Js�W�a��sI&rkؚ��9n���2�Y,���4���
7ɳ$j����ٳG�߻��;?�z�o��ʱ#ǧ&&�_�z�����175�N��C��b��V�J���$����/�85�k��R[�6o������m��ٙ9kD��)y#y�����lÌ��p�jԄCU`1�x�B=U�J=��np���Oc�T��6e��Y�f-���4+�Z�i������
G~���ǐ�Z��pJ��S~ ��nZ�W��4tя�32�N�f�;U��ӭ�4z�"C͊��{)i�a�+���%��{����4<�(Æ*r�ܶD���)1���'��Е�VS[M�&�P:qH�r�¨ך|
���)��a�2�$���/����!�q륥�۷oCW�}�[PI���[֮]s쟘l|�{�;}�%�������ow���z��s����c^=�^��V�J9�'
�	�i��׾V��8�i�R@`�!���W�2�p��撰��j��n ��3W���=_��B@��Y�F���_ɓ�fg������$J]�m�3+�|k�5ױ ! ��pP��f�6j��~��^�b}D�8R �ą*f�i��������2ʒl �)��/�B\{�e ��\�rk�:�<X�O� �xI�K��VGQ�@�D��P����"c� `��D=+�[�^˫�����F��8/�(L�(jifz�u-�T� S��T?�\�b�A�녶{.������
�[/KM�JE��Բ!�Pj�6:�t��VQ�S�l$lZb�{+�uJ��hYյ:��Z:��d!�����t\�~���_)֫�b�!�D�H�.G#c���O�Ih�B���D2�Q��0����d�^(MPN4��1�C��55D-� s�|��p"$/Na\�q*""��2��U�t�W��}X*���v$���c��CI��WWY����0�Ub�L�h���,	=^�����1H\�9��ɓ'�cS��z��!gaF�x޿���:u�&����,xexX�x�TC"&gø�z�*>�߿�w����w��Xrx��Ǐ�4Z���c<��k���xF�E����j3��xpR2����:i�Z?=z����>���E��կ~E���v��#HJ��.����;w���1	��"0����&>��A���񈅧X1�ٹ����ͯߜ��931~���K�Gf�n��Ti�Σ��Aݨz�͍��� ��j��G��O nk��g���{v����S��+�Ն�8�4��&�6�u�����v���A۲�4�<w�3cu�f��j��s��u��ᇌ�h�]M��b6L�
yZ><K���l��:��$`��	�m��,�#�8N��jk����	��I`���0*H{��iH�	�	s�N^� ��9�,;�i/��.�M��l��*���Yn��[� ��	߰��p2�CUlr��0Qf�A�*ۑ�K��t=�x���-n��&�M�kn6�:���^9w��׾^kMe=�y��-�[oE'�<p���1י�z�F2�T��$v�헅��Ys�;�<��ZI�n������A�^�v��i_�� <�d]�6Nx1\����s�M��6������L"�7�,X�*G�Tx��ѝD�Mk�:�N H!<�~�mȜ��z�[[*�᭬�� (V�j�:��@�CT�[�i�E��^s��0�掫2'�~����f~�3�F1j�N���̐��gذ��������l?���Zc��VT�����<������À�&s�.t���b��2�H�^�,K��WE?�]!lL�L�.�f�\�U�$�������L�t��~������׿���{�����\��1��(��,x�����K����SRe5{�������^:w��8���L�������	�6,]B\���8��i����/aͿY����Uj�u��I?͓��5cx�c-ᯀ�Z�d�Dj(%�z����=հ
�+MU��r�:_4�87�ܭ۞�hFJ��]`�M��M���B�P��!.U��'�T�(\�����O��$��į��8W�4tw�$T��i^$ʨ�:��?�oD�{��ACH'�1�pr����3�.J�p2���蘌����,�8���V��0�t;�����e��*-�41�X�� *HVE+�k�RF�ti�;��Q��kW�-�o�|�O(�(�UA�S,t�dշ��a1�>|�0��w��JWSl3�DyZ�]Uĥ���[�|�>3�!2�+SY����f4��-�ݻ��Sl��NӘ"F3f:��P�|:�a��	f�~�F��jwmнD/��ׁ�!��p� �Y���o��� q)<���u{�4Ɇ<����d͢�a'rN���h#^�v�
 ����v�E��;�2c���T�xY,�ŭ��4��D��x�=����������"w��$>��!D���s�=(rBG�#줙�p�@0�=����������q/�E���^{��3���^���7�
 �H��boo !/���:C�F��4�%S�:E/#&���w��KV�b˴}K��&W�� ��y�����|���|�+g^\[]���l��\��ݾ�{�3_9�&����#xL�v��*vv���8��1���{*��2�8��������$㊚S^�zՈǳa�j�s���FU��d�K�2��&�i�/�/���O><�"r���Jr:3��%���t=C��6;싘2�2��N�6�?���.�6�3
^�r�1>Y00<W
98?j�K�s�Ej�o�O���B;�&��p���ٓ��kO�wK�V�a�6v�m?�j��K�@�����DG�4�u7��\i����e�H�O���'OV$�˰��4�`΋N:S95[T��
����Π����;췽&���>FP&����k�rE����x�>�oY��x�j�$�8���ݵ�����>�j-��ؽ{�ÇKK+��ݩ��}�����8�i3��$N��B�5F��u�C��m��/hk�&
++}kX|Xt2�ڶ+|��%q�:���d��TaӅ�w�.//C�]�t�������o��뮮.㘅�Ň��y��S�g�}x�[?��h�Q7?]y�sԫ�J[ۮ��g�)G/d5�#`��hRdndI��X
�����lb��ٳ�����H�P^��>0J��MC�%r�����<O,����X����� Tݫ�4�J��E޵�ZxLǋ���r�Ck���:v�h��W�\������w������@�O�� B��b�Py8jBU%�'*#�Ȭ�!�\��:�avo��ݻwC;������b��%���<Y��9.���F;M�����z+8��ss��6�&��8���k�e&a_����N���[�i��w�FoÒH�%Qf&��`r�nڹ ����!*t��v���Ȁ<���`� �u߉-�g�XvaJ��Bm�P���[5��:㼄4�'�fM��S�	�k��[��(s�kO�	��xF��¯���F0+	�(��CNDC�
۠7a�OZ�R�����F��5&dt��垙��tힽ�f��� ��d�N���{�3��hUE�,�^:�J�r��"��D@Y֐���nײ�5Ƿ��7p�����L0y�a��F�V��^K�^l*�������f����][Z}*�q#a��dPڭH�J�B{�q'Ƞ#G��;w�&��6�e,�n�,�~�N�j���8~�Z�a�.�a�n
C�}0�:C�IP�lX�Ȣܝ�$��6A@�Kٍc�����K}���.  a;H7\��_�*	щ��Eئ �����p@&� l�����8���Dld�gϞ����c�+��pkO���_�ȵ7�x���H����4L��&&n��+�0z$���:������Z�� �ݷ��m< T/����?������xF�+���r��eV��,�W��x��ML~�*N�rƋ`��ʘ:#a�bEX��w�n�p;��+K��N��ԩS����+0<6~ŐΜ9�/IAN�$4�A@f�Ji��WI5�w���uU��Ŏ�<G�؋��p�R�;6�n�J�OrG�κ��'�'��yYd��2%}���(���7H�q�8{�f�����`vz�5&fӾ���A|����~��LL�-�<�� B@���z����2
�~�݊e��D}m�1�{ezRZEA�2����G�&n�i���`*�%-A������Ya�rS���KVR�1\C@����s�V�3^7�"�м���i���m������ژ�f}�r:�~b�:	�P��TUhn�p*=)U$Pes�M�Qr�|�8�L����x��_�k�TZ!��XU�[1J'�T�|[�U~n��l�̄vYD?�_nİ❴�%���B�š��Å�F�V�	���ﶓdfbkH�>��@�ޛ^��i$�ߖ���,�,�~����ȓ�HUwq2LJ����MKu5��x؂��Q�(
}u��M�{5I��c�\��ZP�@n��Ҝ�Lp����Z�0�~�q��6켴�8L�L��m{����{�oݜ�?v��t!��Ix$��L�O߼qu�L�;`��x�2�C���8��[v��XΒAͭea���di�jM�ͤIy���ɱ�t6�;�=�t_<v�P͎����{�P$
ߨ{>�zwSҳ�u-)���*���c�mAW�s-U���i����������z�׿y{yiѷM�㭍���x )2�lT�}�X����,�H�L����N��;�A8?Y{R�Տ?�r\���C�V��̳���i�ǩ^4��ƺ��
��RY{�*h:4uȴ�t�A����Y�(��N���x�w�ą��>�����I������ٹgzrjjl�s����\������ONN�L��üV\�v�H��p5���[;v��b!ɐ繰� !�<�?�VK�h̨�]_5t�i�z�
���c��˩��s/�{�������+�����=s��A\���P��Ò�����%��A~��Uqe���%< fuuu0ȓ42K��"��n��� }`$��	��'�cqӳf!��a�ُ����8����m����������������3j�D3�<�\�BJc�G�0ɣ�Բ(����:L�^�	099f����9�h�C�
�ͺ뉶��\:B�`��5  #����q��ў�q�BU�ؖj���\��"[NJ>q�IU�@�6ؒ\�P�eGa��>�ų�:e������n�Eh�N�!�B�����m+o7���S�Cxv>3�� �-���ݕuq*�^%:ֱ�<��O�����$
O ������2�cv�G�ߟ�c�iE���S���� �y���S��lc�6��~rzB�11]g���� ����K0�1X�0�0*�g���,曑þڣ@Kg�%:��Ρj^;�p�9��Ma�SsC�0�J��ZX#D���~He����������2~�r�
�`����p�r�{0, �Zy�9`\w�4qK��E ]�� �Ih���:�6�����W���/
�sW� LL��|�EJtɬ)�I'��)@/��2����0�y�<�׿�������
n���j�������qY`�00��",����Z�s� �%G�5 D��HZ k O�Ka������cF.K���̟?��+���I&�2;����J�}/^$\g��f ���
�`I�i�N����T�������n�X$���W�5����JTN��=y����5�Nw�5��m,��|//$ι����Q����[�������3�ñ}gqy%�>x���g���aXF��E ��0� ������>PeWr�L�)LbI(RZ�y���X�CX�w4}裭r=�2AyX�Ҋ5uUt�)x:�,����b���:�)�n0���%{��3�t�}Co���� ���*�8�V��^�_Fk%�d9��ɣ����uҲL�(��H�t�0�д����c�ԭ�%*m�^ez2�u��4��ؔ����`Nw�!��Pڐ��0����pSQ��P���3Y6���rT<�1ɘU�Dn
����5�r�<-E��~kC����Br�$/U�Kh��&C��5,�,U�&;K�!�)v�!�a-=z���xzI�����G+�K��*C�����@�{A��N�޷w�Ɋ]��J���1�[q�~G@U	L�܈,IQ����h�!��Nw��`���s;� Bf=|d�ֈw\?�˗/C��F��;��$���+l��9�ƻ���۷�����7��M�%f�EIE7�_�����e4?���-�B&wƢU_��Ç�Ζ�������[�yjF�*�݂�x\��s:����n���g��5#�.�1F��t+�j�0��m�m��:F=����A��u�ر����k�?��1W���ǋ��#������ݼ{Gj�[�j,�q��%\�ԩ�9r�X��b�q���铀�}t�	u�S�ְ���
� ���R��X���U͡l�,�����ݻ���[���M1;�d����YXXy���T-�Y�m �"-4?���KnT�̈́OU��
����4̕v[��c����qj�ܻgW���az��Un�gy/�-Eɇ|���w���Z����FI�@f����/���j� �m��J_�[,�!}{���R�c
�vƽ�v�iON��+�IXCu�iԂܒP`��/�8I�?�K)h�nU ��J���)��*��i(�nl2�z�9Y��`=`�K,E�"�Ԏ�a�?��L�<�m���Ʊ��R
@�<\�V%}!\�V��ܦ-�O"	~-({lbJA���ˏ?y��������F!�$A��ti#2gk
m��8%#�r �4r���̚�`|���%>K�lo˽Q�b���-q�r���֨�B���M���H���5Ȕ� ��OКW!ӑ�j5'e%%#��x}��a�B(�˂y#�2�:��$�c������ZL�v3>��@A�ba~1Ս��g�,:
24T{�39�F����⎯��*3s��`R�z�MY���btC�b׿��p��VBl�H����	IO<���f:5|���q/|��Zx���F�+ ���7n� z�P�;�+��	���B���	M�8�{�_��xp�[�^���dU�~���۷C���/����ݻǆq|_l�z��\��ld��{c#�(	 �1ux#�j���z뭷t�_k���`,�5q<�sB8�j�/���
P������=��TΞ=�0`�4������/��Q2��z�N�Β�χ+䭮��}�o*Vt(�Mv!1��w�5~���"��;��s�-[f���X����X�����m�{�h97�\$�b��ceT�=iѦz�);�.}��V����70�֘*S�s��V�[�K�JTQ'yՄ]iM�0��B�ш"��:3�e�������'O�d�_� �DD����
�g���cF�)�TDl*חj��r�
z^$'�C|��1k�o=�0 �j�����VPi�R�$�a�`��R�q&O-U�f:��V�y�V�Z�|�Y�o�Ǥ'���a�*b�I��\�N��;*�P!S���Fn[����䶸��>��y��H��K�� �lnَ��.ϋ7�6��)�FZ�oJM=��,�[)�OU�(J�<B�̸�0a.�ܾr9�����,N���
4���0�޼��=W�Y�i�"�,Dhf�����6��ne�06ha�y�?f	��"��#�ҴL¤����/LHŹ}�S�IG���X���P3��Ј���{�^�ьӢ,�ߍ%d�v�U4�ڐ~�\��deuvf��[����?�����'�5�T۟��Ze�qj��
�Y>���� ��/���B���[�o�Y�r
6��&�R���s���,���x��p��T��Q��j��j�m�$�]�[%�҈Q�~��Ec�mpHDSa���I�;�߱s������ R2��/
s��K=���T�x����{�?~���}�CB���J|�-X�Fd���M�`P��`��2}B�����{nu;ׯ�Pw�n�0��]U�t�֭G���ՠ͡(ً\9�J�������2�,��q���eB?J�+-H�RZ�<Ě���E���5������Toszu�ɥK�_~��~�xi��CM6�5ORm��m�pijzǗ��!�䇡	��f��� |�E�u���Nw �xrr|nvrjl6
��k�YW�fa��!stG�8��R�h���l�ͦ�n��Y�+�{$V��YZ��4R����ERg<�l��$VΒ���
� ��A��lda��O��Y�¬X�5I�K1�8K��|��t�������ʓ������`�H3L�&&4�2B�췦"	�`]׆��4Zq6` ) U`I!�Ԥhӂ�ۜ:BB:�~�;��Kg��\z�"
�6��S5orb��7/-P#�t|��4�Ad;|�0 [Y����I�lV]/��0x�������d�s��	Jla�}׮]���7��ܹs�����y�,&�m���$�f|Z��i��S'C�x6O$�������G� op�#������X���l�	�(�%X8�;^Y��#xv��l���k����E�v��	c;M!fW�H83�	��b��a��*\��;lM���,�t��7�$[����m6YA�|�<��/����o~S��a-�s�� p0�����:t<
����܂�Ʉp�}10\�'?�	S�L�����I6�r��Ub>;�hcb�++�pS �����HvQz=Y�D�
�>:��x�i7�l�21p1�HJ��o+�)��� B�����qUt�j4����sH(��N�&��F���m+ˡPW��F��>v�Q^��Rmɇ��7''vi�����'P;П�_��7H��!pҠ���r�ܖ(bi�&ƕ��IwH,�KF�q�Ѧ�2P\6���cn���v;�f�gi S�p�r2$��)�!��$�:�L��Ga-�;wkk �e�YL&=��f?[Ů���ëaC���gh�LN`�Mҁ�*8R����H�>�B	��sX���SJg�0�?m@J$gt����sGrk^���
EX�`kH�o�n�6Ԁ��u�*��(k�@�� ���5�w��\�%����ځ.�lߴp5�5�.H�QMG���7C�/�T4о�n�~���Q͘���� �у�v��!��=�TocXVq�j�#h6�y0���AGyi�Q�fR��&q�<���`R{�ʄ��Q�s��B�e��b\-�W��4Wz���l�rJi�Ǧ�n�6G�ӓ�����q[�+�KX�G`���tG%�)�7����*"44������ʍ�?~�:�4���{p��U�d�0 �4��t{����Y)�})F�����D�ѭΆ�<v�%ԉ���2�:�Q��N��t�URMM����jקvX���2�LYg�W�U�ƚ�`L[�"B�IjR
�Z��z��������98�k�����G�g�1���c�E֜��l܈�1�'�\��+W���?�Pjbb��@V��8�zJ�g�il?�$��As��j<c�:�5�o���[��ߋ�D���[Ѡ��j����b���4�J5ɅN�1R�x��VA��������'썆E���	ct=�epm	 ���"K˩ɉ�/��	���=Y���a����͎����Rs	4�	�/��s�P��@ՙ'�+����)-;�lO%��~�S��n�M6�Y���O>���ʭ[�4�kM���v?�p�1���3���ZC���N%o[Q�aWI���L���$jj�f�J��Z�f���nX��&�M�y�u��(��AB�D�2�l+��o�|��������9�Y,)��
��a~^R��~j�頲k;Jr	�D��	ݛ�f� %F���0���Vѳ,�&;���<Â-�ku)�������\Z넊b�%/"��Ƙ8q٢	o`.�fr�͛7�S�U��[�5d�-,���,j:٩�c�	�זb���;l)(H
X�̃b�>e�����و�~kz+uq��E&*c^d#*�x@�������qk���`X��li�
(�2z���c��ʸ&��ӧOC��p|���L�����ߺu��ѣ���ŋL{ ���!�����I��&�Y�@'�b."[��@���"b\R?44O�<��� 7���)�/q�gp)bHX���G�l����w�]MY)�#?��cߓ+�k���xj���ݻ1��.]�8q �h�y�o�	�r�Lb0�#�v���F:ݾ}��?�)Pܞ={`�����?��_|0	G���;�CVb�.��Q�4��R�rX��6��ILQ������ݹK(�|�rTm"�'-#�R�O?�����nv��$S	����3�����oߞ�p,��i&��U~.�a��[��_1�9��_)�����X�������ɡ���9�f���w��e��&p �O��|-�h<>�ר�qZ�mbh�'����)>�n�AsQ�OgϞ�b�k%
b�+uqƋ��]>�14Q�N��%T��Б�X{D�d��j�?�j��z�����J#��猲ڤ����Rm���ʹeeC�O��� ll/�sXL�`�m6m��|E�L��H��k����0�|2S�Ϸ�8�XI�|���pX>>)TlY��r�#Sz��|25K�n;aw�.�,��pf�V�2rB;L�9��)F�ΨY�t��м�2l`�V���wg���8v\��E�����J��Q��J�
�'�,��1�%� x�(m����JS� �C�b# ��� �ä1V`k�2��ܒ3oJ���cn����fONOM���&q#�`����}!��]ZBJ�ɞRT����V�k[���85Q.5�<��Mi�M��J�.� ��rI���{fvn��ҥ��;���[���Ȅ�P{@�-zt]m��U7��aX&��˦���賠�9ZT�U�CE V�]�Fֲ�n��X�ʆ0����PA+�;w����2&�CA�A$+Jbb��͍�0��A]o����?�裷�y[$�?�b#���i���g��.5PT�H�Ӄ��{�piu�V��������Ǳwi[���[]]Xx$� �5�ʕ6|��\~l\�*��|T�bЎ�y��X����o^f4�5�x�������S�;r�56!����������L4�K�� c!�B�i��m��zP�)<55i'݁���,/.>����n4�b`��?���_ݸpc�	̄�`΀�[Y2�9t�	)��>�C Y���L"�jg�*p�"W�İ�Ke��ح�UOS/L��5��&R)� ���H�����`�XJE$!$9�֩7��:��x��d��1l��J{��
��|�C%*�Mhl��m//���(��u�;���ɴ�~�8L��v���\<$�ڷ��ۧ�h��r��NF����1�"��
����ѣG8���0���X?�ǥhj�E���O������T�b�Ok�(�W#�(�'�造�M)�!�PaCz�΃���8��ޅ�㾀*N�v�	K��?Ý�=lt���;���ЋAy�Ib3�\Ϙ4�K<���49����{������&���a00���י��6���(���1\�Ν;L�}qͯ}�k��?��?c*~��_aV�Ձ��N��_oܸ�S������W�^�~�:C�=�׎�������~�,F̃��m�Yڷo�>@�H����.\x�Wpk��>��)j�wRy���6ᥗ^�T
L����#1r��kB���1��5�#��W��U��>���u54�	e�,��-�FN	&~xۅ� ӆ~�R���3-mM�՟t��e�z�)<�1tŨ��p��?�O��²����������������#���0u⭇���C�J��D��S^�'Q!&�)��?y&�ё}�O�B�%%ku��4�~��&�[��؂ExH�0�� �`���*�/�,�\]Ly�T8at��TU�j�#�#^^�VU�Ij;�|h�1��,-�J96 �0	��D{�m���=x@9��c�)�nbl��kJ���u���FK��@��aCA��?�S��v>�$q��C� ��I�lp�,C�M�.�(hK8J��q<y�RՔIWx#��1U��!����!I\(J�6	l��D�m�.�E"D;E����:@Ԇ�am$�@U����2�"�=�DU��#6V��YV��E�#KmԷ�$S�)��XW
Q�ZbK�M�f{¯y����nd�'66��,y�)8��R7<r��86��q�BO;Y*�޾T��xx�cG��bxm)�5bCel�T�
\��zP�j����f��e^�I���Z�Ն;��Y������Au�wT$�;7H$'N����1LP���-韛`�vJ;��=�!�X��&
SSs��B���?�d)ėbl�ApAb��P-�ˬJgǵT�ճ�㰭E�nK@C�2vHl�2��I��M�a�Rܙ��,���խf9,�V���{��e�w�N�sŊq���r��`a�Y&!"�U��tB���!�-�ȦB.I����ʚ�-���9/�۰`X�<Q��[�%�W��i^�veSq��L�(�5I�M���3>'m�iz,��?W��v��N�-E�8=I�q�:���Y���o�
�r��0�K�D��6���a;���s��S�sػ8i��/���d�J���|Z�U.l���)�i����G��nԏr���y�߈O޺w�ҽ��	�S~1ȒRҍkvY�Cj2��L%.����Bu��8�2I�����$���0{�0F. �G�ip[��&e�B�f���ć#�(�w��iq����R9����s�r�$Y���J�'�Z��f?����-UA(!W���i�y5B�m���H���5�O֒�F,�t�l��#��i<�R�v$�F9�x)�,��N���tvb��F���{�V���*;�f�Ӿ!1K�a�uZ�1��%T���]� ��M�tt�Le���F{�(�)�uoV���>q�4.�Hپ{��e߬H�7$ݗ*XU=F��S�æ����`�~�E�+�l0r��^{�M?�D��`Za~�p �>��M�^x��TpA�3	K�kqq0	��L�a���G�[���)8��6@Gl��-����#�	V,[O��F����s r��ҕZxRi���P�y�x}t��~�;�9y�${�_�1�y�o��&�4�,�`�
�����lL�$� u$$�$	,��'�`~Ht��$^"���$+�+c�o�:��j�N�g��$����,��0!��8�\s�&�������?�#˙��d�Èb9̕<?�L�n�B�E0��7�n��k���dGE%� ��\\�0Q{���AbIi��Kj��Օ��v�Hb���dZPZA�ƙ!V��5�0���I�S�zI�!�w�)$�`�/	Ui�̌����e�!�2
�p������s�|������u{�a҅K�T�fDg�������?d-��5I�C�\��d�e�v]̇�Y�zX�ضݭ@��vd���>���i�]c�w��=��B7	��e��QWD�rK!�OdC/�b�dFH�$�A�llK���jUh�졄�ɶ����$Qi桄B�y����e��АUJ�C�ԕ��fj���Ý0*[܋rMYE�6�5?O�"��Y�vV�F���[ڊQ��Y����R��
=K�l������� ê&%\�\�i�7ƨ���J�(la�q΄���1����`C�A[�^��q�V.�X�=��:Ô�Iϙ�/�ĕ$� �q)�9t23�6��re�9�K\TR�u�|����xs~n@8������pt��dF��������^�;$9�]��)3Y�M`ؘ�8Wt�rX�����ɳ�� d���
w��/0�,��$�>�_�D�w �*�QoCz�������Īii�1_G�tb�Q՝H7%=P���C�zO�}$j��E���̓�S��cI�z���}���wn߄�ؽg���4v,���I�A����DnX6%Ú�xn޾��5����4��:������={˙� �p������
MqX(ǽ�(�eH�j4��FhQ�ZM����K�8NQw`&�Q4�y��tH�h�K#Q��Qy��	V#�Uk�-
ʋ�4(�� SvZb�B��K�.��잞ۻ�v33s_b��&K��[M��
��Se3;x��kw�ޅ� �Bϲ�8�$��b��Ĺ���Z�9���%���\S�
�Lz� ~�g
���h��1Tf�$��G�,���� ~��A"`m)���%��$�an'cG�ϋ\����Ei�ǕU4Hus��4�pw��T��9vz�g�6���	}��j�P�lY�9
�5��h[�)���16�(!"3������So�!h:b����:�c#���<z�H ���i��.�8{�`��(�u:Dji�گx�.\��0�h�ӣϐ�I���m�C��鐆H�`��z��sj��"�fh����+�IJ�q$C�oZ<��㽈��1�ӛR,X�9��%��Y��%��G]�v�1
�g��+� ���10��^�'������{��h� VWWqw<%2;PJo8�C�����W^y��ٳl%A/ �,�7��c�p5��ѩ+��\.
�ކ�B� �a>ϝ;Ǚg<���^�|��������Y�t��yv���M�J��`G)f׮]���pA��ku�R ~0cD��( �8����g܂��EY<�>1����t� �20W>�_�YȾ���RX�-���j�_�G�L���e��f+����)0�+�XF(��:=1<�Բ}j(�v
��P}�d�#���鰋=�,*`�O�ڳ�1�����-��Ir��Q5��(��=,[�q�M(,�f.���Z�|���b,�С4L�j@ӅU����6H����BeKb�+�'3!g�Z�����f���)ȉ^t�㓜O�®
b�`aaG0yR�\:U��0��J
'R��7�2����)�A�x�Su,u�X��f�$,/�r�ߵ��fgk�̬f���eX����YAAìc�`OQ�j��T�3u
&��B�C7��J�he^����\+4%R��;UI�8B�5��0��#���ы���
�|�+�B�Y�~ׇ�O���Q����j�a�u�ՙ��T�t�4���i���\�f~�Q�
<�mTO�#����B,����YiQ�����"߈Vhw�xY���xc�������}kfb�oB~� w�T��`��HҬ�[�ra�-�8�#IE�S�y�^rR���R���4
{ll<IB�w�B��Mz�3s�:t�x�F�-U��nܺ}���{��f�m�N���]]Y�鿓:V������y�'�)l`C)�Bkd��\u�~�˲<&`��ΨC�Iɩ��MtĪMب�{�G��u��6j�,C���W������w���nQ3DC,��H>��)�0l(gJx��b��)�����͛7������d��6$�!��I��=���8�'oApa�bd�*�4�}�Hj\�c��T���a;�Z"{L1w��54551�۔6�Ä��`TҪ�_���2�v=�O6�3Y��b�Β�O�erl<�.9�761s��~Ġ:4���od�ν��:�׾/q�B� B�a��@R:j;~��hy�F-	Z�3NQ��]NXF��5+�f����x�܉�A"�nff�i���MVI�]&�|�mb���O��%S�LUJ<�GRn>�}�ԲBk��b�i+R��G�+	�C���'�#+Mq�9e�z��^F��R۪"ת-]�(�ÀȎtݭNS�M���&8MКk��|���I��PZ�I*�IO���av8��3��]g׃B�f�����M�+I5��Do�-D=�4�2���QRԽZP�5�-h���JVZ�J�������@�.��b��<��X���k-�v��`�3c�ɠ(&�G(�I���`��I(cܰ�aĐI��N�aZ0�9��q�01�5ٔN�! ��G����7��������C<#K� ~��A��=�c`A6�/6B��`b>z�|���
� t ��'}뭷0��֔��.��#;�� ��ظ8cA�@�����1��ϸ�&�H��f�؁�bf�'��AX��w<;y�{�=����� �ů�k�Z�=.c0�㗜l��1Wd;����a�I�eEk���G��&�Lt/��,���)���F"�a�<���
�N0T�� ��1���p &����5dy�&8�M�b��p]X]�/�����׏�~A��jMۭei��gv����}����:Ϩ�p7��FH��kR��2�X^<�����ʚW�d���Y0�QXB���+���ھGN��ޡ"5��&.Lf��J�@�B�a��}�]Eqa�`�2��?莏M�'��C�ڱ[������?i�86L�Le�x�_{���D\*����D���O�~��1o�|�	��Y�B>�mNV��Dw��HE�j�VBL�:u����X������?�f%�\p#Hn�~�{��u,����K�)K}�k��RbaJ��c=-��GyT
�;>5�`�̤E�5�i^���Ti�����ȓ����B�/M��,w�Ԉ��R1"�(��<�53h���2���v$�Z��a=v%�a8V�V��V�����&v���bL������'|��<�%��q5�h;Y�yhA�u���rS���(LL��E���:~�;�����ٰ�^oes=Ks�SA��LRx)O�$Mq�=�">�z���^~��wחW�Y�M�z[[+ݵ��A��p����������@o���=9� ��~�)�������5$��4��^/JPR�v:N����q�p�@~#JB�s�
+�ݭC���w�����6L���:���0���XN��C����:�K/E�����j�_(�(�<)§2c�I鏓����`�(c|�*��t#�w�A
q�R@%�rzz�{3h��s4�����Rg�hk^�
�P��ٱuΛ�7��]Љ���*�0���|t�P��Ս�	�t>����X|<lN���u�RN�n�c�"���@(�T�<�N�\����l�U2�\1�ċ4�صZ�XmA�-"��M�A�=R�*KU}�5e�SY�O���]���������S�]L��7�O�ĄeX�W�`���	�Q����!�T���i��ظ����¢.�+��:|��̬�m�o�B���h�ے!�9���w`��������v�F{�51	��`�s��me3SӰ�`�8t�����_��!�t}N��	Epܦ�e�Y��a���mz�_�%.�0�i�Hs�zG��9���>)��ԋ�ɫ�_�a}�Hv1'-5>�"�GO�p$��� M3��������T�Hv5Ti��6��sq��b7��prY�!J�5>6>U��S���ϙ��l��[�2�7Ö���Ř]V۔�5��j~��L7{T#Ì�ES�o�݆�;67,��w�y@��f���WK����HSmҿBz:��J}���
0�Ỹgg:�,`�4�6x��F
�j������"aē�if���eif�Ҩ�`���|�2[L2?��t�T�l<���`6N��^'�&Y��I�����(���ϟp��QL�>Ɉi�C�������d�xM	l\�٨)>����{�&ˮ�L����9��9+3�*k.�P�� �$��(JJ�u��V;�?�#���C?�����~Q���Aj���H�H̨B�yȪ��;�����͍�AK���D�瞳�>{���5|�\�+	�T.u6�ŋ�R̔c9o��g�g�	M̒������­�𻴧a�x�bZxi\�_�P��v�px�޽+W���7�I�Gl%E J��`H����$端��Oq�`���S��0������(�5�H� ��z�H�n��K�i�4�v	i0�j�~{��)�JV�yen�<2�Z�4D��"�����R��Q6����XY ��º����$��R�i5f0�Ҕ�K!�6��L����ri;>�q�I�	��)(tɯ�#&�a�
��t�f��"M�H��/��(b k�XGt��Ӂ�Ο��E鄟X*X�~����G�p����ǘ�K�|�	�6�����*��mv:s�㹻�v�~d���_d�F+tfV)U1C���$^{��r���7�_<4��YQ�-�3<��L�Dԓe~��$��QɌ'Lr�N=�YI��;��c�;��8�J%�H�:� B��Y/K%�Hm�]�`+�����\��dm��Õ�{�4�*�����8[���9z����������ѽ{�q��q�����K��kK�<�qv����N�<S���K,css[�Qv��nS���BF�H-^i��b������i�[;{w���{������7o��N�k�v���cڮS.��De~z6�]��Zy��bQg�f��J�_�5�w�j���#�ء�ɋ3��ҡ%�&Ƨ�}�c�`
L�����7iZ�^�"w������n��v���+[\�atEi*6R�0��Y�qF��!g�͎��	�8B�$r��l��ǣ5]����t7d� ���:�N��jJ�"��i��X5TL��N(;�G�ΰ8d;�"�i$c��99��"OB��99�����H�N'Ʌ�������༗��57L19P�j�,�<Gq��z"\�p�m�z�2)'` ��0EBG��`�*ঘ;�y�8��lǅ���Tj'OǅH�%䄒d@����x��b�F���V���De]IT(F$�oh�n��{�S�ά���7������G�+���z�ribb|�ة_ ��S�S���LU)�t~����hX�>@N{�	,�f�T��`���_'7bs�&�`�=)k2-�2�vT��c�3굧�W�50+��%z<�Rk���M"w$}��|TM��Y��"���Vj�r��=��q��o���ïj)�w��\kogO���_^�}�1����2HS[�"\K���%٩�y����h^���}�JA�=55�����h2�t���
�0�����?qX�SP��2���UL�5��yQ�9;;��C�Ax���� Z��|��w��!���vr�ţT$Eow�y܁�GBr �h�=����$]1e�1�D�c��S�$CV��<��դp�)D�ǒPf&��l�l���&��HE}[�+��
�N-�h�	���QE7hrB��	�Iժi�8!�3f>��FϺza����y����d��I�@n�{�ON�L�X<d��9��D����=���4��l��\�~`IXw��3,�'������8�ϗ�Ï�\nff�U.�ͩ����<�@P��s�C!7���%��>㄁�q��lÊ�e�0�z^i&]�F0&�	W�")W��%��ӡV�EݜJ��৥���j�z�z��)�*v%�}w�M��K�X�U.I�D\�Xqy�����)΃gJH?*��a�a�(��䀳\w�T�.c���.^��3�T�'�k���I�?��_|��l���u�o��8b�S��\̌���p��a�-�c�����{���!\k�a�H;��@w��t%��x����Zml���~�[-���}�������S(��th�I*�H�,&U���U�ژ�Ҳ���͔����Qo�f��sa+�kC�N�Z�RI����d�I;�T{����2����^g}e�����_{u�T[�[(W+~�<53=��0y��fTnz��������X��kO��~w�٘R����uZ�f�\Y[Y��^�����^?�t���q���)eW���b�se�݅���a�ǚ�c�N�F���k;Bk�ػ�w�~���w����[�U�J춅�kw���� ��z���H��(���.c�ðc8�n��U��"k�/
����᧟>w���x�%U����WW�ed��&�N��z�d�ɥT�?M�SL���^�ȌF y���~��������ql�^����Uh���UR���6�Z"�	q�BYǒK���S�<:�s�M| kN�]th�.]�[�������P�c�򧨭�%ЙNĐV#�cs78,#���#zQ)��j!/���5����{׽u�[�ZM5�O�Q�k�K� ?����j�C�]��V���\��W}�ş�zeW8܋���K8�M���[�Ȼ��	XS�R^*�;=�s�+[V�o�L�#�NS�g��ʤKX����[��&E���;�{м����~�ٙſ�(�7�x���߽}�\£0f��^��+�z��>A���7I��RD�"�-GzMga�Ӵ��Yj�������Y����q�T�!��4�hfs�����X��Q� ;@Ŀ;䁐"��dYE���"r�� ���Pt��S.3uC�߮0��V�G��rU���BA�>X�9T�֔#0m��a�8���i��ք�!���=�P������#�(3�:ʄL�1�O�ٸ%h�c���}�6Cx��=Ǐ���O~�(B��-͚l]�.eb��>M�&�l��ZXX�`�HbO��J�{0� Ѯ��h��7YC/�t0G�����of�Z��fL���r���`[�"��	���fm�?K�a7����,#!ڧ�eE)�
�,cDĮ�e�(u�s�����en���J$7g�>��I#�+��VZ:��W���$G�l�åB�A��B:�q���$��G�_a~p�Re�_�6���'�677G��L/�$Y"���X$З�m�ql�3.0!���O<݈]�@.�V-��7[l������Pc�c������\
�Q-�A�����|J�*&��d�0�?�1'5E��4�'��$�5�}�%�0�V�&���l���O�8~���4��TQ\�eP�6TP?VؾJf�ZMr,qؑ#GN�8A�8|[����|ooGqI�Oz7�0��$�U>�g�y�ܹs�T�N�t ���b~�Q��hpB���Z]���t�i):���A��>LF����C�����1c;�XO�^��-,*�����2�����^g���yz��˿��gOg�M�oqa�fy�K���)�t��M�8r_�Z�î�1��NK.�e��mvو�5I����&�Ͱ����&f��rĕ�	+s��n�	<2��2K��G�Pk�ԩ��^{��J�R�HQ�it�&g^�����?��Ʀ�Zi����$7fg������"w{s�I��`�D�Tz�5������[���f`�o߾P\+��Eh�'�r�)|	������Օ��굱A������>��SF���W>�|���XW�F5;�=���u�봙P�F���s�҉S��f��*vٷ�����sn��>H�`����*B�"m�c��9
��n[�~��e�~L�g�-��n�P�H2/�Mf��'\H�tJr�I�}nO�K@�u�Ç�U�j�R�����w)�Xs�m��,6�@�HO{��PW�QS���0��O<Pk��H���!� ?�>����q����Xf~�!��>Em8�^���HڈLE��UGRf$1�o[u�����bM]K���=�9!���4���*�<�<-�>�v(jh{dy��Uol�rK�4��m�έ5�~�>e���"��9�m'�%�1�j�9}Ju��R%I���m�@Ƿߏ�R.S��\�vυq����JPM�Ҽ���(;3<|�0�[7�>\�kאָ��=B՛o�����MM��vv�7��-;~�\��)$型`�gz%���5I2m����!�Ru�m�X�i�u�,4,Õȋ���f�x�W�*�23 bI���\l&�mz`�w�~Q��Ȓ$"�I�Ҷ�GYߋ4 o�(�
�����؎� Qb�I�Pb�٧N����V!]�G!ˌ&߫�á��\%�(+�4�(�5��!��2aK�s��*p�Aq����an��e��Z&��?o޼y�Ν�zaK����5���]Z]� ]h�	<t�$&)/>�Y�9X*��cX�DA�M����Gh��O'���+�4�ѓO���3t)Q��a)P1Q�O��d�G��0"��ώ`��BM�#�)��"��Ίd����)ˇ8u�I�.�%B ���Z��a�f@�������ΖT��Q�$�SB�"�	�����D�7��@�Mם�A��X)WSi���U��`ձ��1և�0 4���PU7 %0#��x�t9���Q�l
���u�OW�!213I�@:�bW�Z0r��=�l$�p\*r-��M��`�j��y��A�a��;56=1��/~���Z��z3HJ���<H5��*�$�v|���)e�>��s�*r�Ɣց�X2DM����B�@�^�p�F�30���~*nI�8[y�R2p-Z9��O>���f����2!�����:E��R����]��!5�qT.�a��� �T�a��ױ<0x�i�����n�5I��x�Z��0���ۑ �V��R�J��o[F�Qe�,�afjr}c���<|���/?{h�a��Q���1��\�L����h���ʶ��nBQm��Ef =d�w;�pq,�oDF�O���MaTj~9�B
h����@@l���Kf��N��;TL���y��c�;խk׳���`����˶oW'jv����?�����Й�9�|ϰ>����z��w�_�>33��n򒃔g:.�Z��� II�A���'�x �� ���8~hb����A���3�m��z���4��Ź���rk��x�ݷ.]�����z��4���/����������&�<��'�xD#�:�A�Qk���K�|row���yuu�l�����GWW��y�������d�9���+u����P%Rvj��UV�/͇�v���9���}m#� ؎�������˿��K/�4=5�|U��u�[;0\�P9(�dv:�����
 ��t8jt��*)�����]��ah�KT�t*Z1Q�h��fЊR�����@��SuN��Ǡњ>?O^�p0����h&''���^gcm�ݷde*]�{��ĮǮS��{�������:3����Y��p }stk�l1/�w���H�-r�/f��~Fh <,غxj�եʤU'L�\��9@ʞE�tZ��e�')f��ؐ�c��wt��3�j�&4ڞ�����k���������y\<�T��2^ �r��n��1d��Yݶ�!熔�w�{�b^�r
��7Ǫ�W��l��^�sB���Χ�.�S2�4z�ܔ&	�$H�Է��`�*?��,�f��$��u�J��r��h�;���'��[�M2�����w(V�k�
�E��_�E �H�!R��S,-#V��rE��:��0�vw0�$5�E�Rݲ�v���o���w��w���Q��P3��C!l���E��Q���`m�����7i-IO$k�k)�:�^��
Ȕ2/�K�r �r_�OOXa���0+��06��H���N/��_1��@XL�H'-Apeͳ�_�0X���	��$��L�EH`�7qӕܴ��fQ�s�l!0�Y,ԡ�O��v��� B�����A�9�YS/��e��ֹNޣ�|���I��ӭc���HG@��pEzY��c�#���QiN��vw?х�C"�$V2D�T	�0��I� ���Rh��Iݹ�dSLգ�ǐHs�sT���ig�G�u����0l�Eb�G���'�S=q0��Dn�����>��ʎ��x��ǳ��An�L��ԋ�k��26�W`��9S�O�
L|�\U�o�V�!<B)���"�E��ѥ��smeeeg/���$�GP��k�yV4e���,��k`kkGa�
�g*A�bKU&H��������cǎڎ$;v�z��I,T�޵k׸l�>�^���w�إQ'���?��s؞}��;��e�I��LN���Txݸ�@������[��&�şc�16��F��a�R�P�3�TePKi� �VH�^��]ۚ�l�h���cfC�$�W>,�?��o�O>y�С��xc#�����̉�ܒnr��͵̦��d�a����\[[�N�>{r��!�+';ݻWna�sgO����iԪ���Z}�l��ݽ��?�S4�x�.�ۉ�p���p�;u�X�:�>nB�6F�-�^&������{�õ-ǂ&�Ҋ�@�ٙ���C���������Zm�����'���������~���ȗ���!��Z]Yf:JZ1�Ro���R"u�)a�8(u�{�{����`�����Ƶ���͗���N)(��j�V��\߼���l���3Ǐ_����ݍ�j&d)Mc�����u7g�gvw�Q�Dq��ٓ���56�?����ի�d�c�����o��W����27�ٚ�%
��b@\ ���/Z�6u�T�K"j��!�����F1�ڌ�F��������`i��/~�g�Y\8R���`��ݽ{�ƍ��b_�V�� �r�+5�T�|fz�ȑ#KK�>�6$��<�&7��fH�(�{�P�Ou�x�@��b�m��`$�Bos���ՋE��/�z]����˗/�vUR���u)�6��67��^�|Bljz���+ y:�-��J�Q��Ǐ�{�d��۷?���W_}���G�k�cQj����D���4�ܔP�>r�p���^G9�QnǆJb��n?�3�vҒ��k��"G����KS��2��x�5??7ެ9v�޽{XT����"2�A?l�u�8c�q�.�N��扛(�^QA[���P����z-VJ��C D
��NӉ���7o� n�����i7��r��G농A7ʀ'S�b��'��~yz���y��nh�QP�y���w`�5�5f�)󌒗5?�j�@�S��aER�霫�s��Tǂ����`����yz��Hگ�g���f�tZ�����kۏֆ�a7�^JV1��o��>�R��~W̲��H�ז�V�O�B[DX�?��4��-VeVUĆ�t5Q�Hc4�5-Q�	
~���tA�@U��B�� ���Q�΁�b���@�|J�	!KE�X��v2�4(]>����nvQ��)�ŗ^6�בl��h�sy���S�
�3LD�*�MZ��0F�D2Ƃ�a�-WַЬ�m�o�������"
��)�T���%������R��%ׄB�~[qJd�Nd?���#��KE���1��[��M68��Rѡ։.l%�gc(<bhw��	�#�.�q��pߧ;*�!��t�'Ědg��C�HD
]e$�3쎵�LYd�{di�Ȋ,�S�Hi���8�%����VBnP���䂷H�Q�7���������m��bi�(���䳅�9#?����b:�HBM��4�xnV��? O����q&�c¯]��#�����]���ҥ�e<SX$gΜ�z뭷�P�����e� ��v	0;d���8��pK�C�w0�d쵵����M1^G$,r�̽���%���f���֯���`ؔX���'��I�ݽ�����b��kf�1�,g�DD'�'X�����Vn�<K��۷o^~���˘՝�lk�����7+_��?��i�d~3�VVo�4���cA���ٺ��o\��ʾS��/|��g/8�֠��u��lО��ٱ��Yۺ~e�;�땙���4w9R��XSP�F8t;ɦSi�f��#K�]�2�`��?�A��O�7�����a� ].]��l��*}�tEu
w�9�Ε�a��%S�(��}?�������7?��z��G�v�����2<��G��g!��?�ۿ�ϛ��?��Z8̦&�j�zl$Q"D��n\�S��_J���?z�����������ܡc����|�+��n����=��ܼ�@u���c�B���?��_Da_g"�¨%���� -ۢ~g�v1�����8	-[��@�L'NH�b`Xf'O��TjJ��ls|�ܹ��{��ŋT=X̔�X{�����#O�>A*��G�>y��f��.�xj�QW�\Q]�"&��~�"���P'��ޏ�pZ�T��?Ŏ����]ѩ���������Z��0F\�����(_IR*,9�LUS�U� ��8v�4~�`'ǟO?�4���+ѓ�s14�7+Q�&�L��K���0B�><&<2&`�Y��Aa
�gN?YoNR��Z{���uv�����%�����?~�2�5�.���9�t��S�1v�b���6���|��fTd��Ţ��&��IK�%�I;���VMXs]��$��/�ƶ��d��W�>�`ssS5z��#�e�߾}g���;����(ָ�B�Q���<���5���6��9��k�N�<^�B�RZs�J�7�-ϲš��#�@�%����*�ȥ�;���������+������]�4�@����(�6y�Ղ��5R����F�����@��^�T�}ݾ���w��{���n��3>�hd4���T�`�}�f*��� �H�C%zCRH=��Ǥ#&�9��+\wd����<@�b±{!b0?lS���!���	�?�d)�4(&��E���Y*�+�>�0�C�p�m��Ԅa,S�����4�{~���@���:	�.����?��0T/�D2I` ̝��0ā�����V�v���DM;�'��r�S��fq̜zI��z=|��S>�.k�٢���͛�.~7�{z�u&��0QxL�`d	~�q�N	����o�0a]�ڐt8[	a�hn��W#}�H�c�L0�'��,y��K� #i,)�=\�z��4��Q>�'�<=�~#!C��������Q/���p�ɧ������V�����S�=a�aAш��0!�ʞ�H�@�a(��� $%,3e^�
��@	v�a�$����>P0�9�]�A#���BUIF���!������ W_{��H�[&Ƨ0ɷn�Z[[ǐ��U����Κ�3LIϭ�	:��5;;��/\�z��x
 ��붹�(+�Y<a�=�Yu�L��TԮe����X��?س���e	04MN1���Tr��P@��t��ۙd��ٓ��z������w�}��~�~�7~�:5e���O=q����޵˷��Y���Bun��zV�e��2�ex�3ZY�p��ց��<fa�PXv��=S��Jn�����۴����Zm��df��lg}η������K����Rs�J�xg͉�A�x�٠�~������([_{���5ZK�Z`5,�z��ز�rS���Tw�{�ή]���(I����Nsb�W^�s�����/���T��'�,�Lj��~��f�>��L�(hU�������\���>�}}rV�gk�c��?���߿��ڛ�ma���l������{'3ҹ���2v�;�t��w�.�{������͇�+��?���?�5ZJJ�F�@mӉ��z�k���������8��$��m�}�K/P�A4�Z6�>�	�T�S.�b������P�s77� ���F��� Bj[�����~ii	Ҍáa�1�sR��?���7^a�oIM�\B�s����������*��NU�)�:�Mg��/y��Gt1����!Db�.�-�
�2�Y����,����ȷJz�7���_��_ei�\c2�"�F/��>�׋/��2�1�Lx�L��bڟy晥� ֍}�i2�/|���:�b?1�p�,8<��{������2�� �x4���P�y�i<����P�w���G�� �O?�Qouę��ݸu�������&KH����1"d9��E.����c��xD���9i���������0�aӃ��[��`~� ǳ�`�;�e�M�@��S��_��w��A��F/�|4$�}���x��d�-,��x�@%�� r�����?��T��<��uku�� ,;�_A7�Nj����vwk}��K�3���թ�q�Jl+�]`Ӳj=Ո����. ��^we�_���)�Ng� �4�9�w�f�1�B������� �Z+U'0����νFm�V�"�S��1rU��A�*�^�ӓ��F��	r3�ւ*܉���%�����Ky+����#3�g՟=v�������6��ؗ~����I�!+3��h_F��,>��}"��YR��ĉ����^�96��0��R-·��Vh�B5�B�}L�`�>E��N��	i�8X����_�۝hue;��vzߔ�X�f�w������Z�{X�0t`1`��`f�0_��}-ڊD��:pG?����I�N�����t�0�Tc4��)3�Ha���{a�?�.}���03G� PC��4�s�α�7��x��rE�1z�/B&b6���~�i]�M�9|{��7��P��u�)/G�m�D0��}6E��p���<����z�-Ƒ �`q>������{��3�J��+_�
,u|����``��̺���-vq�184F���r����a<��m�1xL` n�;���>����կb�*��׮]#>)z"q�C�DQ���?�я�'��na��t������䓘@Ȳ��~ϝ��g񱒖_���h��
�+��U����ȣv' ��\����GZmH�3Ԫ�'5�Q�Hז4�s#�;Y*U 4�{���z�i*�0ص�WU������$DP�s<��ݲ'�s&Q���f{���Ǫ����*!8�m{(�	��!�����5��I�Nwa���V��k�v�  5u�T/�d��#�,"��j@a�v�޽������˺�Ǝ�-]"E��!F������FTy�L���?�0�.����q�Λ?�	]�Y�NMH�
�e8�6�#H��QN�h�
�����B㣦�্*:J��t;�8q������.���w�@7�9�8���05K����B\�p?γ$�KT#�}o��+1�j�+������ӧ������!6~z��/D��λ��^��Z\�[�Z�-{5���妕���%�$a<��wƺc�>q��47��nqs���'�=q���;{'��i�:Y6���z��Us��!��Q�����cf�۬U�'�kT�\��u���&^z�'g��Nm�������yf�I�Ќ��\�U�n�ݼvgzџ=4�*�����M�ښh@l��~�46��p�|�`���l�q})Y�S�T���=��vK��l�<tݡ�vH3#�� �k@,a3=������-#[Y����k#�����N4��T/r��2������U#wváPN��J��l���qIq���_}sc�l����rc��tw�a�a1�'����e�%�~9^�1&:�F>��f���9�h��G��9�И(OM�di�h3�P55a3�34[� �އ@n"E�V��qj�ԭ��}7��6�^����0�%����R�"	H�f������O/x��r���s�/.���;F��d����l7��gϞ��w�K�}T��U�.f�h2�|�]��hZ�*̝�l�z��.�P`�U?�t���H�'�#��?Ww׏�=vz����Ċ=�N���Ƃw�T�]:v���d(����M�'}����gl5������7���+�j���u ,Uv�o����F����_���d�$�%.ZAO=5���/��R%BΡ���Ƙ�}��'p�N�:Fd���wv׳<�t�YV�Vl򳂖y$I"&]���Lԍ���řT3��N�=rd�T�<XYY_�������چ]RT�8����H�ڨ�I:�@�R��y��rd:��m]���mj��ݸv���/�^�`vv
�����\��k������%����A�W��4��۫�YF}cu����;���B�о]���I]%�IP�z[�9�ܒT0`4���t}o�����Zͯ.dD��I�\<��`��)a��qo;��I67=U�V�����K+~�wqh7��/��Ey,mۓ��%;9���e�d�����`�R�,�9U���n�0��`̹�`:"`@
 �f�ꖅ5�ę*'H�u�5VV�����ؗ^z��6v�˥�֓�;}�Q�F��0	�q,�dMr;$#���L��3����/Ҩ䢭Bl�8��Aa%o��~�5�?:v{�>��t�$u ce�ʌ~X�,naZ�*�')D�b�Y��-��YXL6c�>���2���ZA5�0t!&CvL����;]�Y�Ơ�K�|��6�0v���DsN`� ��Mv8���"+�E[��Q��� �3�O���>M8t�����/������yp�S�N�W_}���o���(�"����������K/;v���w��
p�U�D���-ttIB�j�	g����]*�i��m�S����Ae􆌂D8�7'�Y\\�A�1��!�k�;\"��a$���+��[�=zD~9R&�'q��l(�j�m�7:,�����b�|Y�q��)��(�H�f�1�yz��t1�
�bu�$�OėkO��`v��y�ٓ2�QU�e
F�F^1����i?oFP����+�F��ܩ�7�Ĩ��R������$AP�V���<�����KU�ͪ�PJ�˽v�ȱ�P�wob:om��`#�����u�J���ɶ���~9����1`VЇ���S�/_�$�.�=K����p
��~�:U�J6�h�s1�+�h�i�yny������ŋ���˗/�`l���Sda��IB-�DNf9w����;q��鳺�v���j�{�7�Z-��ӹ��9Q��N�F����� �\\��<����R��*�9b)�z������&`����)����4�j�	<��3",��ߐ�*�y/���i5�c���S����u,�����D�)�%�zn6f��8�(����lT�=J�6>NjJ�i�J��b��<��{�;7�^ XieF��S;��M��v~j�=n����v6%K%��l]�u����dx�F�пQ'I�nkf�>2z���`�R8���R�z|���q��)aO�e��ۖz��`�v7��p�����4�ڐ�x A_(�<kH������c�<�����4n?;4�PU�<1���K��xv����󧦈�{53��J�P�QEx����
�ٰ̔���
l���L��F.�|tsaz��uk
n��ڪc;Z���I�変y�F��.���,�77kc��Tlp����޾u�z�Y����~�ӳ1m���Sذ�TҳbP��+UfhLQ@�VƎ�'s(yt�35]�?T����h"I�;M�B�̒H�X���%�Y�?wX���2P$f��P��#Ȯ�Օ�P�`а��������:dn1��:�9���P���2�B�ۆ
����=�ml�RAj������Օͻw�޹sgyy�t��aY-騇^�Ǖ����h��$?C���B�,���M�/�$���VV����ղ{��I�>�y!њ�#��$(v������n\q��(�\Ӳ�ϴ��6=����J�w�,N�;�p�ԕ���V;#�6O���B�=����s5^i�a��Fҏ���. ��}�*��=WmiID�-��P�~�>�����䂯����I@���qr43f��$�2���Sޅs��}p��Fo��4�NL �ʌ��0<�^��ӓ* �`I	0�.x �v�~�����2�� {��E�sf;�:���M"
�}E�7�y�D{ ���=��K�%�pt��}��P�b	14�I9Y$Ö/�c)?�����4��i�2�1����\�mll��+;�,����H�t���{�� n��p~�
'��!�'0� B����,��w����m6�>�{�C�t�>=s���`�����w��y�T�(�W�y����a�b6��.�}�ٯ~���q��{@,�$>b`��$n
��	���=�dLfl�Ǽ�E����ϋ?�Z>��#�zjV]�C�qV�`$���#!�3Ի4 �Pd��4/�״f�EP�7�Ҋ-�biG�	C��\��A�����&���^�9�h�窯�"P�fb\�ZҤQ)cG���7�q��w*;p'�a�����'7 ���������c�Fj�J�vKq��I�?쏸:���>|���ݱ���:�> g��;�;Y�KN#YZ:z���v��G7wvv��w���X�dN�Fl�_b�qC��;�OO�~�n5&��9{���3��߽v�r���֭�a��dI��bĄc~VV�O���~)�,����|N��!�	�����d�	��N_��-�G�_�0��S'O=�$��0��w\3���n�1m@�յ�Ѱ땍r���j�$�sޒ��0�*u�֬U�^���ѕ�����_*S�4�`ƪ�on��Q�3�Mi�
D��+a��us�21%�c��yɴ�a�@5z�W�K�8�{뾻^ujf�61��9��pE{*�`���;��%���11]�ȓ8,y�s�Y�ꔚ�k�t����4���K^	��Z���N��ʝ^g���$�h�7(���v���و��'N<x�|���a8��a$<׳������,1)`t�6���`�
3K�t��6�	ْ0^�zŖ�[�+��]�5h*�O��k�s�'�.��f�61U�qcww����J����z3VW����Ԇ$����gg���Q�@�N;���'YАP&�j�DWɌ�u	�,MNCb
Ih�p���,��d���r��(���)$�P�ẸY��;E���*}�Z�Cfh?�ֳ�(�%CA�cS�S�xB���\�1bA��<�l�*�U�b̉--ԡ\>BIN#���~+���Cg�J;�v��[�\�Dz�(����o��������ǏC������4����$}���$8i@�w�N��7o���ſ��Wa����qfuGM�~�����n����hdɹ8}r��m��0��+��l�{�0���eB�� 2�L����w���8"aq&�+��	6Q�Y���s���/L~G�;=�	����l��	����3c�Y������F77ׇ��SN�!to�Q���6�o�y��_��׿���k���/"d:�BP�
��7������Y
ܽ~�:��5�%��|a��d �c5��%��V7�<�-h}wjv�B͍j��N�%Ng:�Zk8Hz���JKJ���J
p.�Y@sR[��%���v�V�2�lhB�OV��@a��H�5�92�L��(��%��
9��ʕf�זWzvtd�b�#C_���Y%������@�<�ˈq�}o-���d�j�D�"�`������Ȓ���ۆ���J��V��g#�=vq��q�y�E����E��/?]���jް �8�bx�ǰ��E��D&��i��ED8�i��/JC�A�����(
�{0E�)�3����σ�2�p���Щ�[�����C& Z��lz͖��Ĝ=�/~�����^�v_T�	����*>��sϱv��	ӸY�8ϸ:���=/��2��p�N�߅�ąs���L����Ϛ�r
�N�W�a�G�`~�ҍ��2�f��|��M��u�G��~��
M/AP��mn�t�R��ݥDYj�X &�����
x���#Eq�wL�t�5LMM^D��i��I�~��9��R�^1�Rr�k��M���!���\+%����?���3��߼T��#�e����4P�>	
!T��k��.X�Y����O���o�t��>ns1�w�vy��_|�EL�k���I��+����]8�	��(:��A�0Ӊ�}4�D|��'�����}�]� υHO�ui�Ċ:bG!�ԠX�����r����D��;�ؔw��ȧ�_0-jq%àĞ�B�`��S��[��Pb]�w'��xj]?��M `#w�0������h���B��V�~P�T_o[�Aj��t���i�Ҥld��8;}�������O�P qb�A���J���z8i�sHv�������ͽz�Js�ΥDzw7T�~�p���Xs�W�����ߋS�_�����H@\�pm��.�b�������{��Չ��0	���x�r��.L�R�Fj1z���As�ǁB�Qmb����}y�t��<��O���s����hcm���^��d��	�rF���.^~�K�[���Y����b�Z*k]r�"���jN���l�Ç��ʑ�|��+�j�;�-��G���T)��4���0O�Z�2En�	�ܽ{��!��󩧞�|�	uձ���?��=��n�tq�?��#%�Vˁ/��b����cD�����Fga1MK70
���L��tSuV�Ь/��}¯Q E�`�Ή���׺Q�.�)fd�0N7�&5I��v` E�o����Z�Jj8w��gWKՁ�D)`��Yԃ����j�k�%�2s۔�U\È�����%�:��R���	�QA֑��-���X��a0
W�5=����_��/	�L��>���Ѫ�>x�'o��>d3\e��0�}3)[$�Z��ڊ�:�y������mx�٪�����݇�����I}�b+��FR�c�A�@Z����e�<#%j��}�@�%��v�k{{w �r��H�m�I����*���gnגk{�@ .ES,��+���R��huu�p\H�ϧ��� �+|Evm�\��b�F��:�DiHC�:��V�r��&�������96u$>Cq�ڪ����V�Fj�I�v�+� W�*��\�I�,�S�����	�cK��-4�	]neQ�X��~)�1��E�ڟI�,2���H2���S23� CR�%Y���x�&��Tjv�~��n�=�ϕ�Y��|(HI����Rg�{���4s{}�#�{�iS�ֈT*�~VM�e����j<枊t�v�+��@Q��0��4�`���<�R�{���k��t�@�YO�B��nm��� !-�� um%�:䍡mGiE:i��yg?�~X�D�t^���%�&�a�P����4	l�C��<GR,��MO7g����ce$��0+�}�	�����W�^Ũ`�r�D0Xy-��޸q����@b����^���o��s-//s� �|��ɓ��K����x����Lq��#iTxO����L��GG�a6 a	T��k���{7oބA�o��x�6���^��S%�� F�-(�x��Dg�"� ~�``ff��Ç�/_V�@G��h���ε���'%=�V�\�P�1��I�p��$4I�$F�QFӳ@de�<�Q�T:�L�� �A8�0�9Ӡ�4}��)��ѻ�M�F�Qr��?8|�����޿��0I�|ꋏ�~,Ǝ�^و�~Än��)�f�W���=��Xҥ�Wa�>�:��/��g������mO1XQ]y.AodU�mI�2F�����T��YH�8Gу%�0�Ξ=}���+���`8yG�ͩ��l�K�4+n�%?�!��ݩ��?-c>g,��t[ 9kx>n�,~޻wf7�7�C�f�E��J���}A�J�樃Cy��%r ��n�Y����H��SϞW�A���[g��6d>�2��mM�?�����t�uI��y)�&ݲ=eb	�oރ���!pE�v�V���D�R���&J�+��tJ�"�V�;�V�<Y�;>5u�i�����V4������ڌ�ؐ��Le��xf���楋ˍ�Vk�>6V��>>�t*���A�는NQ��о��$6`{�t#|-��n����_����y����D� a�U��$�&��Xy������j���<X��������;Q���{���67qL�z�����@ED��r�R���U�+�З4-�T�UK��@��Eb�Lk��� �=�xAB@=��c���'��4��ٙ�6�rP�!.}7��F*�r3S�4�(E�T�MM4Be�JH*e�^�㣔�G�jD�>���l|F�"#§������@!ݻ�@�/���C�کQ��HyǊ>'�mW�!��Na�a�0î-�2~�4;;{���\*2B�e��	�������ة\9I�aņf���+��,�\��CukAMyʞ�d�'�+t1���=�v��QD���kk�H��=�H�M�g�\�m�Y�6���3�'���k�&W�������ظ{����&�4`U+R}��*~��EB�=i��K88���),MO�����/�-��!�|I���f&��.d0���԰JP��b������JS����b*`��1��IrB��rU!��R�ˆvp]�0�^�����ݘxto%LB'�}���ar�M�6�3H��LJ�]���O��ȶrO�8V$�>���{[k�sSS�+�~?�b�Rv}�I��.ڶ#�ivT��gBI��1� ��vŻ�}fR�j@�A�v�qh�aR��P�qnJ�_�/y��-�"�#G4C��A�R�l�t�Aؗ"�^'\��
�u~�~�B���ĈQP8���n��T�������|���+�	zh�S|��V�2�A�0_V��G�픔�E�⤻�A���I
Y���Iu)�x�x�xi�O�@Zp��H���pLic��&�㑺FS�+|��ð������yU$�,�x2|��@�9� Aƅ��)	���x�;�(�&�b&1O��q6BGZf8xqq�W^!�"g1g�`�YO�'A��!�1$�ɜ9s�w�k��eii�8����.��@ 7@ȿ��_��2`�1h�t��d�3??�^�x�H̆O!� �96��3�reU"�O*9�~�[�z��0R��[�X��į�گa��P%^���r� ;2����J�)��$��l<�����{d#m_�)�0G�w�!z��ցty]>T�D��W�jH�=�����P�Ұ�ZSұ�?�L� �r�����C���j������`u�]�5d+�����b���[���/bX���4N2cp�����������ڠہ�o��&���{n�2��ǳʕ@��"� B��CL>{������P�2۪�Nʀ�eE�'jXn�*LH�`��I�8w��O���|��o u�K0�-v��OJ>T{�O53I�NU�5?�C���M7�"�,Y��q*�u���q�M,0����څ�eFkL��J-Mc�Xp�e#����5�0��4�K"1l�������н���_�Juղ�R�WS�W�.p0{�Nl�﹉U�v箝��ܴ;V�:Nw�k���f�cG�����\�qk��Q/���xw}=��ƃ�əCn�W=¡v�����kz��G_���3�`��6����j����jn�Į�p�I0�T�֒v�Q�2�y;�ۻ��������8y�@�����U!�O���˶q߄��Z���o�y���Tډ����sa[8rz�P�P�J�8IKc��`����?E�i��nwǕD6�������0�-����T��m&UVA	��ֹ�L��͠\�mg������(�2�$t{R8n��@D�{�ߓv���^�� 5K��!w<T��S� �ٵLSM�,7�$oȘ s���jb�}Y�ٶ2s�IbZ��T��#�>�p��%&WC���'���d96dcDT�}5Q�~zZ R9�~>��ez1�����t�	k�)2�R3�t�0���itT��o��o�Ӌ�V���!>)<A�-�ɱ���R�3�u#Š�% p���Ȣ9A��t*>CI���.��0��S͸4�s�h��9B��ӏ>���߆LV��~��Z�s�!���4�.ro��B�$�j����u�������#�7;�ndZy���R���O���fsRh�Lc�*�4�#�ɔ����LϺ�_��Zc�;�K#����K�Z|O��b'y���+i6�Β.�嚨�\�6�E��AUEҦ��YoЇ�����W�Qi�ia%E��Nx����Fxtbq��Њ[ƙ��C�3j���)�J��%��q�S��Ic�E��&���D�n�^.�E�GGY�Z��gZC�᜘�� �\��a ȅ�MJ��N�ْ�P���ݥ�3�f��v qam�+�i��l�2#�=ˇymt�Q�]���~�]���2)��324�󇃸��2���*����V�U�+�<F��Um��*�U}�;r WX�
-�R�!U1��n{�}��`p�����6��^�����X�P�k�q�cTLV��i�P��c�g؝�c��
\��dcxJw�ѹ�Z���f����c�P�G:$�qādIƟkkk�̃�	�79��ZߐI�R�`Ќ�8q���?��/���,q��Fx E d!�Mx���Ug�gA��H�vJ� �O�<IGE�Pկf����l�g���<�^�w1':�Ƽy�M:)kX���X�8��P9{���˗1�3)n��u ��Ͼ����>>"f&�6+�h�R�㮡K0{�o�f����/��<� �	�90��5��`�6�nv�S(���*�1	*UG�zDBp)�S9��7�nw���8����7����Q�m��R'v���ǎ�ˢ�m�lwa�A�@�5k5/�ޘk$����{��s?����~x���≥c��<X������(�on�W$=>�q��H;�~��J2KبRL&S���U�Q�2�b�������7�� ���*��IyZ2&��]�8����=���q���������-��8�����8�Ӿ��VN6�U���W$���G�y�/�^�(�����<N\$���*���`���(�����v��R��~��Q����@������l��,�^������G���2,7�������z�5{�y�¹�_��N��p{;l�ccu��s����n������Ɩo�&f����1`��vcss���$��|�H��vgc�Ѡ��jV�ZM�p��~dH�̄T:�;���;��U鳾���W+���z&iZ�����TS��Ӟ���`{�ҥ��ì�g� �3�\���R��X�z�<)�pU�%-%�l[~���0L�\+�@@�=�a�|5J����U!�73�})�������q���F
.̇���e����(S%\�vȍ˗��ɟ����zCū�<�g�e����J������R� �?�lR�?m{ff�Ա�N{��������¼_���UGI��KUB�����o޼���~��W_������_~�̙3\�Ω�|�`�{��A��D�8#����B���+VkO��W-2�k����1Ex����W�O�����E�T����j���k��N?q�g�~�V�H����woc~>z�ɧup�:�&��2�v+���h��RZ��ST�#U`�v���:^�]�L��z�8�����IOD7��
ȇ�>}�na +��Ra�����W�
8�{����\���t�N(sQth~�'/<����&�?{��Ϯ��|`aq�Y*�����c���ª*JzHo6 �CeG&�����W�I��җ�r�^j����v���s}NUG9Yfb��\�����x��3�G��ԑ�S�k'i�ĸ���Uϯ�UR��U*K������W�UU��&��\�)�$�0-*؍��[~�YIn�^�{�\!S	�jg�5u}3O +�J �.��ʰ%�@�{�Ij%�'®sD:����v�����=��+nW�/9Qh`TQoШz�a��Wi0�d�}��?? V�[�NS����z���N�2_�����(>XL�-��G�(d�`kN:�MM�<}z����N��tŹ"��5��G�9v��c�tho�f�+��u;:�X��bE&����& �wY�����b�д�G_g�	�J�U��ɋ�bI	����&��q6��,�P�ANĢ۷�	�K`���BUM0�a��y�X�l�igp E!S�Y&�;�=��x܀.�% #�:�/�vL�`�����3�p�·�����e�wS��իtyB��I5����4��z�)~J��ĆB@Sy��~خny��D`0�
w�w�޽��o~�+_��|�� �mM���Ǐ�:Ǜ�ΝÄ��C�k,<��!�7cS�.0kظ0~���������0��wF�i!�E�@�Ϡ��tS�[�$�p؁}�#	�X6�`=�tr����N�Q���gI� ��$}�-�B޵���vj�u��ɗ���G�n��=�4��vO<~���s���Y���p[�6��ČZ��c����pu�������`qv|}c�w���^�R*Y82=?u�έ08��A�cĉ⢵�kׅ9�R+�wq�xv�Ξ�w(e=>ޜ�����v�X�XA�.�4���7u,���8�C�r$���o~s������0��c*�55쵭�m��j��13c�ss!A����?=5.όO�Ziw,���r�bu1ډ7�g��Ng�� �aee��WG4Ez�c�uʁO
DW�R�kE�ȃG�  ug{e�n^�����Zɨ�d��
�6y�N7�$�����ǡ�+^�����4���-�?�ܳN�7�����s_y��p8v�(�Uj��S'�dVڪՏ��+uA��O�=������Su6fd��ۛ;��g����ސ����2SUf2��bb1�*���ܡn_*��/���	�9kXWX��],W&2|Le�,q�������ѻ�󇱋'��;��Guzz
SQ03959պs�Ӝh%k}�̍�a�ر��m�dls�Օ5<�N����U*53��gk��I	�-��pz[&��Ν{�sff�=�p�SSS"��?���[�S�Fk����p!P+����?���O�����{p_����#r��6� ������w�nݢ~��q
)?�/��82=�l�~�6��I�.��1׮]��%��P��q_	�����v{'���ׯ_�,� 1'�JX�Ϊ�9j��b(�@b?��>�bh�o�IT�����W�4 Э��ևT�,A�v�Qz³b�"J��|�ͷ�i�O���٦�������Ӯ�k[[��n}��^[]�����j�=0�����|���ʫ�Ac��\��=< ��1�\#:>*��h�G�'f�ϑ���XL��ɱz�U��N�RZ�J%&�RYd!Y�����t��4��(���%0$�eh^��{�>���Y����.]�t�+�0kv0��m5��e�� �X2�+������_bB.���Y�JqD{Wl	���Y#��zR��]*Ik�~O\c���#�ӭ��X�=y!� FΟ;{ha&M�A�T�>���U�G����mR�i��ۖY����������{��\P;d$�4X��,�۬Z�7Jð��4.��;b�n��%�P��f��0��Vc
�]�����z�ڃ�L�����7��[kb	q�d�TF�������N����X2ͪ��R�5Z*e��c�̓�:�;��/}{}�� <�� 	��H��bQ�=�x&��8.'�%vMUʱ˙*����2��'Q�Ğd�q�dI&%Q��
�  b_޾��}����N�M@r�2]�r��z����]���;���g����&*T~�o7��V{�.ʄk�hVj ��q�2ҍn�N��2W�^m����#f��-�^�̷�_-���@���j*{l��7�){appxy�aR��8ذ�D�������-9-(�e;&�_1�6θ�N�9��Un�#�<yO��
L�#0ld�W��@̭����\�ɕ-��γM՟��3��&�jG�~���p2��A���'\�Y�H�����Rn�0_����0Y�v0� �����ι'�bI,..2O7����u8?L�Z�i�oܸ�-ưq*|�;r9|�q�^�#�w��W�r���Ç!� ���@D�
T#����Œ�=��`͍�=��?��xphǽ{��8�w�}��S���da��C�)^����0����gA���$ؗ{���^�u��� �����;|��8 T�x�{�=L"���$0�\��G��ӄ�����3�}©0��4%,�<�'����?�j��%�{d�+��T��QB� -�`��@ �F��ٔ��)���5����V�aD�i7
��T���KSl�y�n��N��z�����sN�|��g>дLyJz�2�F����z�jD�n��C��}�`��_��a�if�<iq����R|3	���^��^,����3���u�8`�d�U*X�v�qr�h�*A�r�F&��0����9�pob���Q�b�~�ԩ|�׷��M�`3�8�|��C��R<Q-�7�D-�1�j���&�F%+,h��X�Y�	���&��9���$V��%Qτ�?��0��uXR��1�Z4� 'ܑ�2����+j�q1ű�fg���o�Ư9~2�2��g���������1��a�znt�b v�ݸ�ԴQ*�$�XѨ�5&����t�<5�o2j�Z[�@$��]Q,�t�a��=zߣʾ��ZQj+�������cs����Ɓn9qj�ӏ||x�Qg��멣#�5gWJj��{��pr��%'Q��� :"-[qr9z�$ܪ�'�U�ցL�v�A��˗1�P��|!�I��-�P�,�l� �E�=�>2ӗ_|啗^�&��Z���X��b�X
���޲lH$���J�9�� �D<�����8��f'N�~�߭nm9���^]Z[+���)�r�wL����;��yn�N ��-O��(���[���파�RZ[w-����^)r�eE��E 
�FaP��9	T�r����Q���� ��!6>�j�[��@S/���v*���j�ץ�W�n'l�,�+X���H��ZBFݺu{�u
d);�8	�U��޽k�O��O��/���Pa�q�(+P�	�a
�N�a�ɜ�l��3����u/ҧ�O���6�9��ߒUң�V�M�eWֹ2 ��N|�.Q~����-y��6������|�K9xd~p�[~��ٷ�9�9����R-�C�=�Mf��566U�
-_oTq�Ye-�dX՘蠕�5à��V����o��v�����}�S����k�np��;vLLN�NL�ٿ��|���02�+��R�^�ӿ��6A!2"�}�e($�V���_��F�����̸e�,�1����yRp���kޞ��O֔�,-B��ył��)F%��Pf��v윺xq����b�R⥵��v}�v����,��K�|��4#��������hl��������Be���xeokumu�b;���޼���*��	tf�!�'����ݍ��K/�X�u���33#���=�Z�Vm�9orz�R�ӂ�o�Vu� ���N�Vø�w; �Y�t¨��Э���N��.F?��(���Zݨ���˞N��e6}�A������Gn��LhT��m"�6FK�]	��!l���b�퓓7g����[�С�i]��ch0O�+8��k!{�H x��
����;!Ei�"����+6(zM	e�Yg&Gv��|�Av�H�4�p�c��Y����Օ�d������ej�S�0{z����#��)�\4RȲT�|R��3+.����,^���o��0�%��ˋAs|1�����M/{�:"���aqZ�=��O���t�"5���W8G:w�t�Z�~�񜺍'9p� |���Z�4����y�fh<&��� ���8`�?C��2�*ǈp�ɓ'�8̠���/~��\=ŀV����q��#��,<23�r��dN��d�W��|�7`��#G�<��#P�<��4�C��y��8�p��q<�W�� k1,d�ٲ��M9��� ����<� ߘ�A����ī?IC"m�Ea ̸�q������<�E�XÅ#mB݆Q(��f���{�Q�T��&�.F �i뜕J�V�eG)eym���ҕ�7��گ��_;��S���"4����j����G�J�O2Ӧ�W����:1���˗�����ַ��6.G��-7+�ς{8z�}�f���E�X�c�踲$�n}���y�_DI�Չ���9�����TY� ��6P̴�� �,v�tK���*�gf��/`��g�gY�Da$|Ϛ!rJ�y1�_� K慍��
$��
�	Z�8�%%�l<��*�Kj�ŕXR��J�ѩ���	�����B�65�
���fI�ԟy�3W��o-z(�~���X�����!W�6�Xu�0�L�Dܲ�"�'l��3�I[�Hn�I�0��uC*��0#����|T��]�n����@G�;)E�(�l��p���ba朂^Hӡn�I��=8<\�(I��6��g���*e Di�YJ���o�Q����Z�C8��k��aP��46�Vo��$hd�L�8��<�Cw����Z��14]5�ﶒ�3:2�on�Zk�Y����|�45�6���1��lי��^]��ʋ߁�+�7�����Oⴄ$�6������"�u,/(��j��8,������T��t-ԍdp�@D�j:>F5���V��C�Tz�27�̊C�l����	-p]+��퐯v-FsʁY��G�g~ �u�����Pe2��8s��[�Z \���5l7�/{9����/�H�@�OC4A��p�0FF��ˍ�a�C�c�ANrȺ��#�ʥ�H�G�cHVI:P��(�vzS/@S���;d7�~~N.���OƓ5�T�!��Ի�Ε-\�
�#�������R6�ֆ����mc��ݘhl ��Ϟ=��_�xj�ĉP�����/�z��N�pz<t4��I�����x�T�T.ZEKKd�4똄ťۿ����[��[�v�Є�౰���%�b�}������O_��_~�)�&��m׵��~+�G�}���b��
v��f���y�S9���3�I[�N���f���T*�i2�u ɮ��x�� u��{&��R��a�N�F�'���@��?�iՖ�3��{��>$���m�:��b�B�+t�v�V��ꄐR�Jw�(�Ag��n}l|qqyii�+�4�+L~T�j܉�&>6�kZZ��Z"k��ū�](�*�QP#ӡ���P�q�.Պm`�V�ȓ��0��Gj�Ti��)Dj>����qc�Vo
��b �6\����ٽ�Ȥ!�].���--�0�2-��g�F�8�+9��5�s�C�=��g�1���ZUa�1w
m�iz�&y/�A��G5���s vz��/z��mB(�*��蟨,V��{;��)�2�h�q\r6����x>�Z�mX�&�$���/��GΤgܯ ��q� �1�1��d�<{�����? ��h���2�g#��e��b`OKF���!�{�k��>e{M��b��~n�I����d�_��kp-N���֟���f7>a�v>�JP���"�̊�h�� � 9 %R��>��+���_F?p�w#�!��w�>��\K0���ݻ�!�s�._�l�I̜&��d���s�9��_\ˌ��˪�c�\Rű��A�_�p���B������kR��9��t�қo�	������m���fp�<�Lw��ٜO�/]�~�����C�nH��<�w�I�l~
���rL�-�b�-:�G�E�(ڶ�Y!�xHyw��#c��
�ʛ��i��0(�3�BN#>+}c�j8�'>z����o|��Ww��P2?�.^��G�>��ʙb�,����˷C(�dp�2=3�V�n/.伒�)�f#���M`,��;�-��sU+�>(�8U�J�I#}ckq~�߉`�-A��;�T(���O���F��W�o����]?�MqT�o����U�[�GiЪ����.�3�D����΅�[m�+
���(�w"M�$lS�p5�}ôe��]9r\��3��}(�rOIk��3�6y�T�����$jW�����o-m|�ɧ���+z��������k+##Cq�ɔedQ�_���Rs�q�����u�ݭe�N��hv}w�42;U,����W���+�;;61|��wy[P��$�����F�4J�l:�PT�C��y�ˢ �&�zjXT�D�����P�
�>D�쓖Fa4��Z�v_!_j�[��G�gwL�^�U�-�(\5��|�%�&?�+��ck�	�!�h�i��ţ�ퟞ�n���)�73�6E��ա�Nld�<v�ŋ��*1%e�����
����B.�ni_��c����;�1�)�DC�Ba� ��;VG���%Q�	C?S� �'|Md��nr��2��R-
Rwۤ D�]��BI&�A�qJp�\f���ֶ��H�ǀ����(����HL�� �����M|�;�ԋ����P2�Fi�Z,��� �9��355�=9I& �W��ȌԿ2�Î$e�q����'7b%�i�S����N����D���_e$�w���΢d�܅ 3,���^�%��3fc�8�N�T ���%�,g'��{�W^/|�!����b����_\\��\�vM�dޠ(�2����K�i�B�k6�������_��_�����Q�
�1�*�l4LaY�2;;������/aZf�w��n.g�>K���G��4=��q��O%�M��SO��o��Q=��#�Bizz�ʕ��[^�5>^�����狺��;��+����g�?��ϏO߸z��܄��LGF��M����`-�P�����7_|�ŷ�:��ې-������]s�6���=�CÎ��!Q���mǱʥ�����`�nX�a�N�°eZ������Y����Mn@�v�3��Ta���M�*"�
6eh�S�sK�ݤ��0Ȉk[�v?��P*�Y�o���}ه��F7`���O=T�*1�hQѫ�6��(rl��T�]n�'O|��Ͷ�2w��aG!Bm;�2ya�#Bdi��ظ�LRA��KcS�F:�HF�	EL۔���t/�F��mǕ}	������{HXf6sK�R"^��u�TI�06��g�˅�###sssKKK7n��Ç��g[�/$�	�(��q�����]YL�����dǎ|��7W�p�0v��Hn�ɢ��*��&COw�9b��������25�S�`��v�V ܓ�b�q0q���7���5���0���;�g��.��Z\$�q0ւ�"�~Hғ'Or4�	��ڹs�x9r��{ܺuo}�Q��������SO=u���>� ��pA�3��LB.�bMɷ�Ӈ{���I�wb,�X��>B&Q��@1�戝z���4��dO�>�_11�$�R�H�(Z�Q����y�#\�)���=k_��'#�R{�"f	Aqf^u@~LK�d��O��t`�'1�0�V��[C#N��L�O�el�o�"����hP��f�������{��w����ғO}��?�lU��6�������+���`�DU5y�uӂ)��Y�v�y�J�U�F�*�`��l7Zd�XZ�>�<���Ij�r�С���R[]]�2 #kɥd)�2��׿�:%6=1)\`�k{t��JbR|�A�P�S�=�es�Ƶ^xC�cn	P� �����I-bb�z�P����S�4WO��V�+bq�B�a��{mƜ.,l&�6��t��X������[�2Kǳ�͔v�M�&(S��7mC�"�R��/?�g���'?�jД��эfcia�����rN�0T��R&g���V�wv�ڼ~�q� �ho^T�C�cy�<����so�������]��>�!����X<���wެ.��=��ɱ�T��_�Z�r�8:T޹��"5����6�G��w����2m�P:��x�ى�a�|��Q�;�v�ƚ��@��z˔�<#���pʞd6]1��C���]'g��|L�qa�6](W��~*y]ɳCN��E.�hX���$�y���%��z��ުmK�O~�ƒ���5,a�i\'^?\������|��^n ������V�A���<L�KׯA��s,L	�^�d�誱�@��R�k(2.qdKP�9i������u$ ⽴�3('�u:z���`!������(s9��񱭞|�IlU���}���vh,`�����9��O����Y@|Q��\6����䒖�r��e�:�`I.�x���ݰ"ഋ~��@Ї�i_�|����z�o�w��%��(�el|xyyekk��)����(�ƨ�W�p�/(�o���H$b;:x�@�R^ZZd?/7�'o��d�Ǆ��q�J���:u�7~�?��b��r�+KD�mY]q��J|�)�0�����W|��o@�A��ޯX�m6Q~���ä�s��l���B�ӫW�c�gg�{����w�;Ӭnݶ����fv�`\y�� ��ɱ�O����7��@�h�bS)c���Ml���=|�qEy�'~򕗾�G����ƫ/u�-=-�׶F�'au��978��rܭo,�1ԇ�CE�zV��&i��dJ?�à�j�ja�H� Q���鄰pw�N#����AaM8�t�W�ȏ�[�!�D���4]�çQP_!���k���KD��%1��i�b%��P܈� )$�=Un�H%;1�.�TB�����F�V7L� J�n��Z*Tza-5��G�X
0^��GFtGi,,�j`@AD��I�f4�Ds�):'��ڐ��d�BDƨ7�d/���B�4!�Ӭ9Ja���"KYxA�A��۷off�U��ڻ�S@[��atı&>?,-����_�?��=قa>�m�
� P �8��d8���B��e�	[XR�{L��e��]������C+N�+2Mn�� �)�����F7==��x��Y_nWʌ�p|$+8�Bw�p�8?Sl�=J��[bj��t���d(�Ç��X&�Ř ���3}�0X��:?�0����}������<1���`L�wqBX����S'�B�|�.I<k�
#N!�H~��L���YU���;8����&�`RZ< ,r��g���᩹�$q8��`j 8�Sa^x�eB�]$��><��8>)[��`��e�F���4��KJ�0z��71�O}���\��RȀ��*'�U�(��&6eL����2��������W�?��ɟ�ɟ2tk�֊��t�w,
�;�N,aZ:0X Xn56�e�fu�VS���\>_,�VoW1 y7��Jk��O��O���	�XH#�1���k�n޸1;;K��(����z�c�S���&VF	3�I��B��� �q1����'?�l��{� aeV���+���XD���(c�M��������&g0�X�^���/^���L�x���W_���0��+]����\�p��T�%Bzg�o���%���Tj'��6�Zl�L�"C͒�Xعc�g?�,.���0:6�Ҟ�^�+���(	�<	}�TS�'�<�R�kk� )"��I7�ۊ�������Nz��|�����,�s��J֗�L�?�X��d��\�`���MÆt����ZP��2�7V�7.��t61�;Pb���g� .��B5 
�I!�P��JM#��8�
�YO��L�Vv��醲�^�,��A���*r�[�kT�*�Ra���}���X�R��6�$�q����V��Uc�L�̧:�:�cΦ�T9�8_�L=U�@���U���[h�0J���G�(�w�$06�}�h���-ǍӨ�n�R,�c9C��)Aק����,m�5�q���8��5�����%�E�� ���ı/x�ʚ�c~~^�;��\�m����W���A��$aDȒ���|��c�@;�r�ڭy !
 RR�E�ի��W9��� �����" e��s;w��e��@��?���Y+qČJ�������)�M����d�PD*P��c�Ƭ2�\ K�=�ѿa�	9��iղ�u?_?O�l������������IhLJR+R\���j�K��]�j�<�G��;�݁�� C��Q*��o3����BhHu�ҩv#I9����_���כ�M�1/_�q��իWӈ�9ÿ2P��$��j`�<��c��ȍ��U�:�GJ;��8'�����t|���~7�m��<�0,�]�5��i|86>��Ё���,n�# !_�U�{M��@V�������=�MG���Wryott�M�B����Kؠ	�C��5�x)��	[�H��.�8L����@%AJ�	�L����Q��Oh��j$���*J���Tj�fB�h�tDB6}���`V"��Q���7ǋv�eKUeI�^�o��sU��V����w*�11$�6�'�+O���iv��]�6S�Q!�:�(��Վ1!�J�o��榝3���� ���-k
�}�}/
���,gMgS.�0.�����@D���6�����@|ܼy�5D0�6�} �fnnB����L������B�H8��yoN���d����&E��M9�ĉL�����A6O`6	�8��K��4�(�Px��IXf8�W�9xd&�`)�1A���qEF2@�ȇ�pţG�rW>�Q��hC����x4|��� �10�5Y�`��o��6�70~��؏�Š��o��Ӟ:u
��gL���i�cp��e���?�t&��Uv�q�ș3gp$�(J�9��ˀu0���a:�?�-�
�}�G05���z�ݖ7n�8~�����p{�H���9�D����ʑeKL�ǀD� �&���(ёT`<�rc�r0Pv3�Bb���j�h�4�}�6,��>�tehв�b��LA��;����0��8�%����!�q��ܵsv|b�������'�ʹ��7ow;q��^Xs-�\�Os���[p���Rik�23R7�n�q��J�:X����${!!�g�}��g�I��n)�VK8���ʞC�$��+�0�*�>���˕F�vj� �,����[1Ss�.��njxC�|�g��S�UL�&gu�F�6�ɏ^*��i62{���S�$��C3{#�i:��܁ ��}Q�}�X������<5<}wH�4U�0��&�h����|�D�4U���%O�QE�����k;�b!��.\�����s?;::N8���Q�G���P*�F��>̢vm֪#�F	��e���R��,�T�m��Yڿ[7��������w�Z�����a���ާ�������C͝viO����76{*������r� �莡W�l�64��#n��Hm��gʨ���jZ��h8��:�K�����p��Sn���t�����\[�{؄6N��i�o�qk�ۺ.Ȃ�eG���,k�#N���m{N����m#����Fscmc3Lc׳Je/�`dF9�.��F�� ���ǟ�7�  �+�37��ŋY���A�_)�\��-��C?&L���ڦcyq���4S!�ۭ6�`�����U]�ME�� lB_����M=��	��a@�"J�Wey!�Xn�هxvsĄ1\,$"���~��v�@i�s�i*D�	�@��>�=�D�����m�kKK+".Q��1��;��	a������ɷ�zeh�D�h�Gf1e���Xc��@����'�ns�;$�YvogU�"1z�|rN7��nw�`�+���,'�3���Keâ�Hb3�@�P�����?���{�:tddd�}d��MN�r'<>��֭[�G�XQ���rz+�I�F��A�v���A葓��3ʭ	'g�~���Sh�(�J�
������ӧ��O�=����TKd���L�8q��Ç��v�OM	G6U���o������/�4?'d�����-($���'j�6�d�������r�n�Q\�j�����oޜ�����ׯh��Sׯ�/�\�`�������F�!ô�V6�/<�Z�2<�Üd``"Z��ô2��
,n��wC��L&����m�;aJk'��̄�����5�_�`�ш_H���=εL� ��.\��D����I�љ�]�.�������z����q���H��r�))���6�j5�f���Z�zf��xȌ>��DD��Zk�����o����zMw�0c�˰(��E�ċ��q;�Oi!��	=�P�C!W�TDKe� �X��)��$��>r�>�	�4����$Ț��q.����J���&�[V��,��pM6qc��a�OMMup�(�*C];v���Kl�s���_X�e1g����f$�$N�%���L��A	�:�+b�.�'�Fр�[P�W|�)�p<n؀�&�ۓel��| ]ȷǼsF|��AN��/���[x�}T������Å�]`��g��ڵ��ß ���9ǒ!�¶;�XY9#:�QZ�J"> �ǓrGI����C+�g�뀆�� ��×_~�;�b�sL$�=�H��M_�6��g!kq�8��X_��`���%;L�L���>�2�_�K��X���]�O�/�ng����-��Q�SE��!�m_�(���ho�3w�A�@�ȀR�n'�@�]�xajv���P���j��j�FۏB�tʃ0��V[�-��� �D��Zv�P4m#L��F���$�k@2q704*�9.
���x���� *�*.W3�A�.�}NN�/�Ҩw��@O��`�Z�-����99��W0�G.�A� �M?0�1E9G�X����f�_)ڎ�l�?�Vm�Т���P�Hj�-�dW;g��UJ������?���%,ٹ���;��v�Uv� ?�IS��x#���D���%0	�Mϱs�Ge��а����o~�;�c�ү�g�b�|�ё7۝<��Y^]m��4�o-l9��j�
���RD��d	���X�s��s�3��5��M!�G�ʠ�d� �V�6��ªm�5h@<)4�����ҍI�֮#�y��|��z���ʆQ���RPtSU�,�'I�fA�ZXh ��n����ek1@���igE�Q(�I�{y7�wU=+�=������R)��ǁF����Zq����J�cC�(���*aJ$ �;~�3�ܷg2��bq&�Jf�� i�[[�w6�R�4=��?t��Wz�q��r���z�����ۙ��3���;jk�G�h3�� ����r�V2JI��V{dn'�g[�n@�[8:΄cBtσܵ����	j�̘�+� H@�������j7訢�<��͛�cc#؇���	�lǳ6a������!��&�K�r�n{aq����P!I�or�����/]�R.9P��\����1��L� o�/�s����9E�����g)������e�,�+/&K��^g�k����d\`g�]���T�~Ro�'���J��������9�k��$�+NQa���3���ɧ� v����g��;\�)ٝ�֟�C�Z-�Z�(#��#'���>��n74��U����Ͽ��k/A�nm^YZZ��v����W0�O}�c��˿|������Gٵs������/�o���Q�%�� ��g��eT&JLͪm{i������f}�ڬ�s�t�Q�99:=^v,�;��=x��޹�~;�ⵝ�+���Z;��ˢ���"J����hotC��u�H4���j�����T| �(��%
>�jL�F��QD�jFQ!��@XHQEj��Pr�3���h��ZVM(3ڐ��C�̓��d�(;�B,�W\��N�P�_S�^�N7�4=�� @�6�C�oW����㺒�s�X�]�4� HY�m�JF�[� �Gp���9�ݕY4�7�r�E��y�:�(b�V�=S��K��
��{^K��ȅ4�[�@&�?�����\��;��2��Y�����8� Y#$�K���<]�������Qh&�	
���{��Vx����������VXQ��6�����6���+�pr6�� -ne�@�1 Ӛ�x������^��`��R��P��o�>��l7�aķN�>��wl�s��o~� B����9x��?��?�_�[�	�M@x�+��9�����/^�ĥq�011��^��pE�<8Άsb���+#R����	C;�g��˒��pN�>��㜸a<2n�{����Ç�}�����w�y��v�Ν��8E����� ��ۘ/#ϭ� �����[��:�g�,s�e�}$�bN��u��Je11��!���c�<p�'ۦ�p����aY����*0��%wdE�5�j�2c���C% ?�jYZ,[���NL�m*b�*�(�LѺa`������H��,��4����5�6�5(4���h>�'"���g�K!i�ϳg�a�LNP/��ׯSZK����$�:��C=%x��ebZ�_�bƚ�F{����!F�RR�<56!��0y4�0�o��=^9�zsbr��qjeH_.������V�ɏ=����[X���������#��ugڨQ	��A:Q��jP�y*����铔�w�y��k���M`c+A9Z:IAⶣ �����Z���j8Llv��6|�r&`�s��+�7sW�{f $0��ʫT%�N�V
�و��E��k�j�kN���_K����륢�:l�V{m)n�d�M)l�Vk��Ak�m�&]#�-ҍ -PD�K<=�`͋RH�8P��rM#U�{rAT�j�F-XZZ�(�\�5�ڐ���o
/��Q�9��N�X"�Xa�(-� HTx�h̡���htB��w�J��Qk7]�y��'�;z��l�;[��ڨөolժ[�i8^H��G�9t�>Mw�(ð�BV�cO=����}��o���.��[v(Ow���I��oU7G��c��;�o��*�Q����n��w�a׶2vuPz*��)Y��x���FCս�W���қ��Q:��m��	����5sWӅ�:ݻ	vƩ,��/��^��L��:n$���=P��{8q�D!ր,���pC9�m�z��	$� bN9��#�bd#��vj2?��HB#i��\hVC�������1�P��f��/)�i���3�g������˙x�b�H>t*�>s�= ������$t�]��Đi�ֈ;JV$��)��w1䣒�{���h�2-J�dΡf��3 ��_��s��{��)8y�NR������z�7(+��񗋷����N�8a�(~�駟�9 ���u���  /�N�=�2�U�~Ёܣ�\�h��z։Z�[�A��I C	�/:�~ �#���?�F��ymemsqycxh��c��''�F��~�B�fjO�)@� 1�A���`�d���6^ɬ���y߶��;�F�&{�Q'�R"�΁{F�J���1�żj�-�吗����� �9�Yz�Z�-�,8�{0���@��V�LھB�p�m�j��;XSq���NF�W��Ut�9d��U3AW銚�Y_�^�ޕө
�mw[K�rWU�n6}��X��Oa�()�l�CL�g�$,d/�ͤ��I�@d�)D����� ����缂�'j�^æ5�u���*�ZӅ�df��ju��ԆO���Ǝ� �����Ё�u#r�#B�� 2U���#�"�_Ɇ�L�Å(�87DU�0''S1.�©`g�W��.������lw���e���-f�U�4s1K#p����y���!ן��m��	�u?s�TB�w�a~�]\1���2�Y�sY.�-�d���V��Ν������z���q ��(fATn,afa|H�:V�xC��≠i�:�3�9q_���z�-�_�U`s&��^���@��?��?���o&1�+l���{�~��_�S�0�<�`Nl{��p�x������_�\3χ�\H"I�Ϡ-G����kt/#��v7`<�E�@�u �<X��~ء�I�*���	y=�4m/�b"'�P5�?�1 M�v�C�=X���rN!���3��QlK�:q��Y�h��r=��b4�76��vH^��[ZY����GGZ^��m�O����:6�R9���'�ʨ�s�w�w�]��o�lڵ�5�\��}�/����זW�#��N�X�N���Fa����o�������ڪ��A3��En@Iٰ��k�������i�:y{�n�ot�"��cof|r�R�`���D���������L����UNǽ��2q�D1g-���FJT��'y�k��Z�ׂ�PB���2t[��V���<�W��Q!���3	�z�Z,UDꓑ#_��h����p1�Wk@#��
~X���j� �����C�n���q�f�����B1�ن�vs^2�g�7��q���R��\����5j+�L�V�>0�Ɲ<��%���$fô��������U(�Vw�.�'w����ߴ���R#��M��Z{+J���VJ
Ł��)3o)[�na�wxHW[A�L�<ӄ�щ���Gʵ�Y/�J0�����4}�_��_߬:��S��xyh4����~Ӱ�(Q�������f�rE`�D44���a�	���?�c�x�c�:��[o��jq��t���j�@��}l��7֖����~���Eu�D��Рi�k!ТI�òMϸ:��*�6:y��{P���_:{n>ގ�@m��rmwڵ�{e���-*M3��"J�rщ+J��Q+!zX.�UE�&��� �?�f)�7ZL�C�"�.7����D�G�A3؛�΁s��m�_�ո��ۑ=|${����ݻh��y�e2C2VF�=�t��s:S(IN�q<��rU�K�Zf&`#��$���6-*�y^\�K������9# ~SH,jrE=R9郳!X����333���c1��O{"E�!�� ���|��@Mr���ٵ͍�ݹ���:-�J�n�ܼu�<P��9�����Z*�%^��.�v>���R����z|zRբLu�G�v��}��{�M��v���h���A���wsE�ݎ\�I���LK�o6����/��i���v6s����{����7��˗������ݿ���Z��ו2�8P`�X�F1�(e_� $�0L�x�:P��0X���ׅ?U�N�;[jD
���`H�3�u���8�F�( �b������i/����2�k�2�7+(o/�E��G� �;�8�ˢ��N[�z�R!�>C�MK�l%i�B�}��ql��"S�}��a/j�a��P���"���'q�&2b=�����r��{Y0�����q&W�s�1+���:���n��G��g׮]�.[�ؼ�p�&$�/�[-9���{��3gdU=L���)|Wd|r��	��B0�l�Q�L��Z�T2~Jo�pw �cfKZ"7�<pT�9ذ�;�,��r#�H�qLI��d�Nf�c���qO!��JbvrV<\�3�Z���c�����g& �K�Wgt*Kce�K�$B�20n	%)����Ǫ+^<h\�ģ��N�? l�Ck��[�
�2�(�D;\��ѣ@J8��ٳg�arr��4qW6��:(bZmf����+L�D��*C�����q���Y�܃�!=w��#��(p͒"�X(U�B���J��i��Bexl|qi��z������q�5���Z�;w�u���pT���V�6I�����o���c�L�#욨�����h����D����^�D�A�X��J�[���+�V�����E+˂��#��羒��g�S�>���+W^}�U���$q��0S�A+�Z���"�I��a�5�*���|�ЛF��X�#�p�z�,-^+�f�P�ȏ�Y<==}j�aX���s��o���k1qt������oܸ27��1q�:6^�c"�V�,'���L��+o'����]z��Ί���\�XS���8����\)���@��q��߼U�7�M�:��F������@� �`Ut)'#�<'�w�Z�̥+�3�Eǌ�a}��|�:����N-W�6r��P~(�DU3�Y9�++�G����Z��N�)�?wV��0�;au����E���q��[5������0�={w��hu}�yv`������ L$kE���k�0�0�!�\�A����Bq��fG�o:^@d��Py��:NDHi�CFg�۱�+�U*���8��������V\Q����q����\�]>����x�P������SQ�,�I�nDO��D�k�6f/�j�Q}j�OL��醣c�a@����}���Ca��������t���f�Ɉ�*��d����w�\�����b����͢˒��̆qc3[���0�̼��c�p�?5�/��d6V�dΰG�G���:�^�gI4����孴%X�J�f����c���溝Iuё�ЋU�h�sA2ƍI����	B)OAW*%`!~:�5�Y�@Q�&��f��{�(�N%Y�CT�sS�O<�9�Z]7W�P��4X[Y�P1��Si;_�2-�o���E.`�pͽ��~$�l1���8?�枽��a%��jvW66��/��mC�Z������{�ڻ���]_���Mځ��Ta+�
%�Z�Ƥ�(:�)���9��Ld}�����%ׄAm�{�)A]�	�ׅ��)�eEA�0���j�0�Sh�Pz�J=JV�Q7��P,���*ѹ����I�Ǒ�i)��UDe�4RӂᢑώL+]����7c�ļ���X(��N��T��G����Y���C	�'�n7��pKv���g�4a3-i��pB/	[���+�e ���+W��ȓ'O�ݻ�ܹs���\N��f ��g1	^���{rTLE4/�,ؐZwʼ����ߟ��;p� S&p�NZ��=v�T�fX�\�"C���_��/*���dJ�,#� ��X�KB^���*n�){,��y��d��l�-�,���.�����b�"(ԟ�,�!xvd����!�xJ�@n�##���,�3�}s���8-Sp['V�|~|�u>�P*�&�x��S�O-���_~��'�|�G�|�!\�?���{��S6��i�<�����C�3<�|K��t��*����\6ǐ�#Zߋi:��%����,�={wc���q<��C8$"�P$a��F]�ɣA؝$�����z�=7{�D9�|�[߁->=�k��}��0��L_o�T�UŰ*#��Ο��� :� ���=<:ގ��o�]?L��]=r���C�QM�YH`*�E��,�,b�M���(�x�;C�����3������Ο?����p�ۮm�-�LL槟��dv�q�Kڵ���$�4P�Z��a�0TX3>� W*�����a����SO���ڭ�������������mvÅ��K��ݚ���E�9���*3;��V�����~k��\�A���}	r�H��E�5�D�p������fsק�]�v</�c��#��][^Z�,�[ZX�r��#�M95\'�]&X����� [ �i��F��L�{�h�yv�E�5m~��J��Y��p��S���ݪ�:݊��F6|f66��_��B ��Հ`��M��aI5��,�p2�����7!ɣ����~g��W�\����G5Mn;�"$���d�G�_��g��ېb�N��0gj~����\)����DY����(=�H��c ]b8�A�&��J���HI7׷�p��
q����&�AA�8LR���6/?�hn��[&f_�t�K�R�5�{��%�Ѱ��N��=���G�+0<�{pp��T9W\�u�H�EeL�_�z/׳\���/%
���P��ߑ�!\n�^k��ر�e�B�Oh+�@����V
%��ON�D;Ĵ����_[���Kb�g�L�	�d�?��Q�C���W�s����]�A'=�����8� �$]�/[����aPFW�p�&�1��Qb������ti��U�0���jZ:���if{y��e*��&+Di��H�`ft���D�Bb�W�^��7�66�>�J��f�I�>�
 �`�h�ئ*�>dMu����(�Wf����$��_�}�����w���X^��w�kW۲�Z�V�� ����5����GB=�t�x�4ov�m�H���Z�:Mq��n4�D��,�,�J���"��z��e���:0��� Q�e�N��P>Y�$�;@6�)�=�"t3�4�ϊV�Z���걜J_�vR֔8y
�S�`2q&��K��ޢ�<s6 �iok�������5JÀ���}r�"eN?bDHҩYT*E~Ti@��
�|�4�:5�R?\k��B05B��F]�^=�l�2t���w/�$B
�Ja��سg���(���W�07��� w&i����A�AX@$ɻ�o�͸B^X$ኯ���zjj
߂!�~|��p�Ç�)`��O8L��e�n���~�9R�?$K�d��,2�a"��1��o�Ɏ.��ª?F!��K���]j�5u��Mb�_#i�ؓ�7Ʀ?_�� �'''9.�����e�6'��0��b���$u�9�>���	لT2\3�6G�x�dr����W�����XKL��þ���1�6O1O�3(b���x|~2�%C=�]���Hۅ�\RI����*���6n��0�˘Ԍ����Fe�9v2%)�8	K�<w����/8z
��Y3�E�ȫ�ejI)��\��ԉOQϼ�.��S�|��C_�x��݄������fff�=�gU���7�h^�T�q�u�ҧ&'����Qԫ�Cʿ���#G��.����������V��h��~��	qW,y��=|����ⵅ�M��f�jh&>��0h��y�mi�g��.OL�=z ������7�Ɖ���w��53�i7�~}����?�g>��_�����O�li�6F)���%J�ɱwe�h��)��h�gEm[��g��}A�%6E� ±t��0�D���T�T�T�4�=
Ň~�J�|K{����sK[�!LQ��~�^BFڡ��*��5�FK�|6]Eu:�j�ury�i�)�Aߴ��F��$j��N}����u�����-e3]������/4G�1�/����tk|�����Qf��1%�s"j��0����y?t`z�V����e�O��2�z�G�WX,�x�\-���{���&�L�����ES�&�������d��M�ԉ��BE��"��n�t�6�����b�jP0F���L�U�o���sg%�ur ��b��I�fa�s�Fm���386Xraeh�v���i�&�Mm�$.T/@�p'�N$2�Dև����4꛼�-ˈ�����c�ڪ��}���Ĉ�����0�"Y	����g?[تV�b�D|�г�v*W�rki�q�� |���8ք5�o�>,�3g�@Pcks��<��.@��Sɬ���齽�d���XG0T`y+ˌ	^<�Iً�դAqy-�{������[6Z��,�s�6����cZ�V�>Oc|>3;�ς�`�����+�
;���R� L%�������P|?���]a;�Lt,B�������w�Qʸ���t r��B��mٰ7�2,�xl�d�/��ؠ�wU�&�mAwc!��%�#��:7��P(a��L�V�Y̹��*�0IZf�t_���GB�P � �Fm@��[tsfA)t��K^!W04űl�n�%�F��k���>�`��]��kq;R%d-+-�� �*�x�r�c��_����v�O֬3l�0M4Y���.�IQ����� ���ȍ��͂�Y����^��^�+U���., ?"����YJ����<,�3�o����Į��A;�%*{�D)�v�z��+w����y�	@�8ĝ����gM۳_෮\���2�Ά ga����i211�`���
a��n���c��,F�!����� ÎMy�he匤��N,�����yxxx��ݸw��a�(a�p��܉'�b�O˥,gϞ=w��a�(H�`���?.,�+�LV�0��E&��rL�d�;u�qx����Q>3_��a=�?t1a�*4{�XpKu"}]8:}�xA�����+hY6��g���c����a`����}�޽���.\�F1"eNDh��ŋ�*KO�-�^7n�*�Y�{Ǐ��o}�&N�x��wށ)�ϹM8;�8!��d����Pd��$g��X��UٴJ�Fes@	��� Cb`�ت`�
L�l��t�6���G�/(�Đ::F�?1=r�ҥo��W�R���G._9����n�햯k������56�f���r��G�����'&:]��i����J�>P���1�Q�ߍ�5�og0�������9�+*q�ln�A�����J43���O|zρ}Ju�ua��\����yO~�X	�[��ǆ>x���ѹ�qغ�����$������86=�Q�m�s��?���n��������''��멧?���ώM�@��۷w}s�m�q����~7v�&?��@�N��L��SrGKC���N ���8Q��������O���*��u���p��7��Μy��'��;72ZP�-���������bd~�Y[Zul�29��Au��R��)"��:D;�G>�8���բ�zG��Vu��@ĭ�|�#^�,��,���˗Οs���CZ��΅˧Ø��32хX7s0��~ӱCP=J��iJ�+<El���uӦ�)�� ��!��)	j�e�1�͋���Y��RJ\b��n���<��jQ�s�V�j�k--�f�W/]>s���R���<ۄ"�*���s���N�9��xeb��w�B��6�9������I�E[}��WN=zbxv���&m���c�Pr�1?O��n�2�ô�/}6(%I'��vZm(y��q<3������ܬJ:�~y��2IΈ�Y��5�����������q�f$@�8O�>��[o���W�U.���_��,;�F�اй��l�BǷn��4gv�DGf�ɒ����T92��5�Jĸ��P�i�K���:��p?��f8�5xe�΀���{xG!�clw�c�S��K�k�O�rj����pQ�˳�f�G��`����v�ۻ�+���������ׯ^�����'��~e�OV�q���?,h�]�r�"{{)��D�[����Ag�Ad`i�*�]s;���,(�oE+ꏨ� L�^v4э�^{�ubrs���;wNc��8-�*C�#�iu�UW﵇�H��m���È�xTr�v;-�5v��~�'
��H�#K�Q���]H�Y�,C�9���+sؽG���=�� '�r���ܶ��h
m��<Q��<=�ltBj�-r�SlN
\�E�b��cZԯ�$01�(Y�T�y��\!�����(�vj��kU�2:[������N���a���E]��Wc(�/�^�9SLb��Flkj�&����n��{9a��.#Ԅ�4x�d��E2��c3��.1�v:gΜ�����2??�ɸ��&���å�l+s@��W��4t�s�%�(�R�|�ԩS�h�2f4��91S�Ը�T���p�7�ޓW�O���HI�&��9GQ��8��5l�� Z�6��IQ?��0�j~vFS����Ird&V6�����Wl�s �������莣�	fffy2M�3�#	��9i8��'~�'�]�������0��|~�P���'<���V��.�'�
�n����
�����5c�X�K:WV�25N����<6$!����dH�*s.��D&��25��i�d�J�]I�5QDݛ��*���´(�������7��ԧ�'FK��w3դ*�|K��ת�ι�xz�v��x�\ιf���9����h�����ݰ�l7U����3M���!����L]׃(�t����3�D�&���?<99]٪��f�4x{q�k_�:6��?�yl1Ζ�K���-��;�'G'!��aT'Y�h'Jb��B;�+Wn��6���#�;w��c\k[����._d>��#��ᱩv�@���ޙ�7�k�f�sTk��g}|������J�^i�����_pWR��#u�*��5��Pa�����~oc}�G�¹p��w���._
���s_�����cw���>�N�uM�w��_j�oM�������Ԑ�a�i��R[_]���]�n���LJ��9#���F5�v*#����i�C�c�� ֊���;���k���XN��԰-�K��(�v��/eDmx��E�'�zr��=��ԣO!�w؍��F�;$۴�[Mܕsȭr�|�R�X����,�;0\��zs�Q��g��ARML���߻t�ͷ\HjЕ���N�4n0��^�r�ڕRe�֍���?x�P��Z�ۢgI�V���7\���Ă���J��?�vCXu�f�K]�D����Wn�J%æ��;v�8p�`� !���Kr3�aKw;a�ձu����.C��B#ro������@�?/3������^��K/��g?;+����Y�%�u%�s���jx��B�
� � 	��`S"�v��+l��!G��?�������և��[2[��y Gb �*T��W��s���g�{�� �;n�|q�޼�'O���^{X�Y�, H{��H|���!�;� Ϝ9�"I&��@�A6-�����f`fFZ�0]�T=����q6��C��C:�}�4�E���
��tV�v-�b?�8�g_w%���j;r�j�l?p�A���LO�ۻ*VYKA�5��1&dB� �%ܔDEɬ�tjzr���w:|�G8r�,~<KH0`��o���ɓ�qe��&m�� c�ɑ"@��0%��ڵkP�R�^H���Q�ًC�=�_��B<�z�dKZF�w�⾽*�*���	)��ۄa�[	�[d]��N���_�����<p����g._>wa��UG	!ؒ���������������نc96+
~�����S_�������ki����&)"��4��d�BV�c�U[菕�#R�0��9^a�L	���]��;�Ҥ����e�>l�a��"���HA'�����tЕ��p 4�e��*CڪT]U���b�onzy>533���mt������+ד�ߘ�LӬմ7�t/>�9�8;�5��?15�R�W:����k���%�kK�x��P��|����nh>��D!3�{�v��b��60���0E��N�>-n`��P����F6j�.pQ�-ӎ�I/�ٱ:�B)L"H����C��{�0���aĀt�L�S�f�[[[X@)�(T$�,'ޠ.��dP�c�>�#�AĮ�cTlÊ�QY�ѐpkՂ��^��=ͧG�I���`��ESp�'��x�s�CfY�.�?��G3��C<�+�E�#�d������WXP0 ����qhb�^\$�yD�@��~D�'M��9�'�a�	SA�:V�Q����V!�BtŚ�ܣ�֔�\ND2|�D��6�����^�pe��%���dy �`����s�Lq��&��4�c��-��� ���j4oܼ���|���*N������]�t�G?���7gw��"�R��]�$"������ji$�ӭAw����5ɟd�))�FݐTUxV
i�b�J��8�?�������jc*���W����_H�J�����]�v-.�u�j)Y��oicjbrvru�ʍ�e����v* �.�
��� �0��b����;4;=_Fy����&3s���կ~�������g`�e��f!�7o�^�v#D�j��4���DZ#��4�l�����(�Ɵ�e�*m-�$�\�GO�����{�'�c��WU�7y��ٯ��dv�\����]����?Z�����_�ܱ�(mL�8^��ШR�MLO�7W�֯��c���<�h@ct�Q���11-�X�Y�m49=	���d�Л��Xܗ�uL�입��q��؃q��`r�?�,�ڞ=F�ЩidZ��Zfea">1iF������݋wNLL�%��R�,@>%4:p�Y�>��WJ�Tf:�?~b��Я��(�~�����a5�|sk=�mY�5g��|wc�{�ݽ{7�Z����%���n;���8ڜ���j����,T|G|�����j3.���f���~sy{���JC��\7UPT��x��temu���h��r)����?t�i�'��؛�g}�K�mg���-�6~��7��4��L� `PG��b{����˘'�-���ܜ�6ǹ�;0 RuIΰ��x�����N�·'N�`�U젝;w��x�>R�IJ�n3�}|�!�m�n�CF]A���6��6�6Q���:[�j��跽�R�膕0=1y����s;w�2��ז���t��\ބ�:~ױ��Ef0[A�~-��=���|��l���gi�+����c�Y�J+B��җ�AhD�d�B4�$���8K��zBX���=Su$�{�fz�9;5��SO��w��E�5aM�O�?	Y¨�R�g�-ʢ�����?��\��+�>�O~�ɵ��O�{��һ뛛�����2���L�c�!(�&[9q�_��������77�/CS�^#
���V�e�U%7х����@D�O*��T�%~k�-FM�eHgV�&y�W�؎�8�c!�L���Ȃ���V4-R�I����v�_a��&�����gLL4�+T��\�XT��hovr���r��U�RUI1��,�"RM`��3SԽI�ۚY�Q65U1�h����)%�0��\q3���2we7&4	n�y�	��: I#�='d�93�4�v$��t����2�Y�������G?
݆�!��Dt��+}cc�@�yVZ�j��B��*R��y��7��}�Q@/\��3S�8f�o\#��E,��X�t��]�"Y�U�.+ܬ���8l�)���ŋ8S�D`0��L�
�B(�P-J��5��z�$n
#��#���1j�Q��L"�6Js*҈�ڟG����O/oG�R�RLU�3�ak� �� �a�gΜ�p�R�j�K�+���0QP�$���g�W)�gMM�<::�4sۘq�wz��a��	�t��f	3�z\褩m�t<�	*�9&�%���ӧΐ0���j �%�Tu��J&7|)l,!���/gϞ}N����.	��S�@gN�<\��N�>��o|�5�hX� J<��t7!��}��Ƒ���罸��&�`�Q! �@��\"N������.,,z[��gs 8I@����9����ȹhí-a���kn`7�ˆ;Y�0�S{ ��L8�W\�[F����J��kMΪ�׶g�I$L�5�:3;_o���� ���3���a���3g��hjr�4\zs�W7�����4���u�è����t�u�.�V��6����Z��������c���g�yN-o�'_X]�61ٺ�{|�#��x��ɦ�svF��R��c(;3�F���gv̸YԪf��5�e�kIm'~����}P�fm6���*]���&��I#N�AX��ٚ��Ne��ѹ�+�j�DQ~m~��G{�+�x;O �{�".}�����^�-Xh�we����Ȣ�TE��� i)��8#w�D��a�4o��@c*/3)��8��o@��p��C[�ޙӧ��8������N�~�K��1=�l�<�����8�� l��U�i�V{�6�8zf�I����gv�]8[^#��X�~�Ĵ����9Ϩ@�z�F����k��N/]��ڛ/F���?��;�Ϊ�[s;f���dsT�l(9����л�a��ϣ�������=�?T�ɧ GU�3�س���c�X�����ٳ�~衇XٯX�,m$��8�������k_c��FGW�ǿ���6jYR������K��8T�}��ُt	c(*G�幎��G�t�n䓟�䗿�{L���^�������?�������?��}��l N��]@P��?*���z�ԧl��\n�[?�s\7Ox/R�N�Y���.�� �^~��Ku)��`�mdud��OL4�9~�N�ڄ���
x�J��v���H#"Q�,��W_�e��?�������K�Wӵu�I���Y$�n/sNMmot��uL�➝��rL1�l���dm���x���.�{��l�hN��~��Fb��s�_�!2��	 �-iK��d���7�HM_����[P���6|'�SK��"}�a6u���Nw+�u)5�R�a�hL9��n����ۉ�`��C�&��ʉW���t�<�R?�nfn �w­�jG����ݻ���q�۪�*�7����!>lAYy��^(rx����U��6!��Gа�פb��m�S�L%�3uD���g:F�XB��-���q�C�i�	]s8��q\�oZ�n��`�򲼄Y�4ԭ^w�x,W���~8Ω����q�`�F�'�'yE)�W�Ν��r�ȑ��Bv�k� �(_�$Ɩ^�\�q���C�������"�>�����u������L�ęx3-���Es?�tf�Ξ={�inܸ�Ӓ�
V>PL"h/bE�� ���<OJ9�.طo��*��,2�&�>�����o�!&�bC$^�s��3���.��M��u�	h5hٹs',��R�_��$�1 >>\��q<Rp$	~����%+��1p�0!�>mbr_�_6�e��q���UX���4�q���$-�©pG�*r��_��r��sE ��9��B�x�����x�,�eL���d��r����Ɇ5��>`j����[���33q��V�����@N�i/W��ZK1�8��-l�f�7c#����*��k��6;9��b�k&"4v�uz��];��u�,�\��U�ΒR�;��*�Jm���:��J�Zs�֥�����gw�e,��a]�[��v���)�èG]ӫT[�啫[k��n\9ph屢�`�Dqǰ�����tR�5lN����صs_s��4UïM��@���[i�f)	r�f�n���oԜ�D�&ao#�3�1���A���A��+7��~w�h������.��<z�����-z%4�G�]�ܕ�rqb)f?C�����	2MWuӌ�g��o�*B��BnI1षw�d/���S�rkȚ����{�����^�q.�~�����$w��*ɚ)�D��$�Μ�s3ZAs�^d*\�)�l����٨Sw�Y(륜�I��R��n�N����\�L���̺� ��R'(\���N�[ɡ<̖[�F˄)5Om�l4aV��~l�I��{�����{Ͽ{5�f� �J�ޜ����N��߻vu	6%p8� ���$��m���E�C�:)��,��D�V����w�������j�������~mϾ=�ɉ��{��z<!��C��
91f�&vr'��V���`r���3L��E����pi �&y_����{� l>I�wma.�d;f�Y��ۘ8t�x�78��;�y��ŷڃt�����A���SG�skk9/�����XI��c�x�#��xօ�CzUWe��T-L�Oɛ�vF$f��#��~��ꇪ��'����%Wf*0l��4�o����n_�W�RZ4���C�))WWvs0�b.��]��;���QB'���Ve>���g�c���	����m	�jq! G@��"n=Fq�	�X)���0�aT�-8=��V��E��N�p�*&f��w�GdM	�k��s��9H��%�����\\0,ӭ�~�95AY��,/H��*�ls���P�߇^cE"�(HO��5B��*��l�a�szQ�J%�4�>tx����y��{Nyߪ�Sǃ�7�,k��j���MU�nA�׋�ucc����u#��?�8{$'ss�.�V�Y`�_}�쵕�������>&��aN�'��1-S�i����W���Þ����L������Z�e�۶L�u�;��}}y}} ��'���� �Vkf���ז��X����������fKk~�r- ��/Q����W"	5�_I���@*X%�;��O�@<A�)i�4�@��\�8�{g�bwv��Zws�n<[8m�4O�����US�(�%��(�ސb�4ʣ.�������܁_Zח�~�Y����y��z�ׇ�«�*�
Uy;�Ɛ�_��@��n���d�Y�1�|�3t�Z�)���1��r�����xb��v�mnn���Vؚ�"�D2:Kh��N� xp�ԩ����5\��%lPF�u����ް����0'�}a_�x������pQX���G��4}13��	!��+��`8q����/�ɠ=r''���ŷlA��n�7��`�?���ᇸ.~u�w�"���0RJ`lO=�>�x�g�~�a|����~���ⴸ
&
�x��J*�RQKKK?��Op_8���(�7�Y�Lf�6	��k�.�D:??�JN����G|$��@|�׻��	R�!�0�#a�q�x��u��i��ߏq��?���g�Wm�/,{�3��O��9�����̙!@�1gϞe��f�&%��n�H0f��@Ά!a،��x&R�~��;��`|ˬB2F�����`���L_��i�Q^:���þk>`��א������Q��`V9q�u}e�򍛝(�D�֥���F?���ȱ�k~k���b�X�S���&�@�
��\�U��@�%f�тA����$�<v���:�ؖ��y�@�	|��ڝ΁Ç������/D�� Q�QJ�D<���vjQ��&pB���P.~��E��BSg���C<�L&�vf^t66W�6<l�V�(77�l˽~���ڲkezLۉf�ȤY%���9��Ĵo�Ő��۽�:<����4B{���rѠg�0G�f�{�ee&� =�,��S�^�t�U�o�.omx����_�S�`r���/Q�<L��k�*���|ū�������%*�M��G����a� U�>���E�(Ff��ET٨g��P�]���Ĥl���5��9V�	&r{*3ìh�ڹ�����?>�����EA���j�Â���:�,��A�%,�2S�ٕ��ۈ���RF+��H��$�bb�ќ�\�t�}����g��c��ȱ�V-K�g����M�+T`h�Z응	|�=�>�g�X:R���T�d*��!�I��L=�B�v��'!o�~h�X}��d�5K���vy�c�UK�p�J':H���ìF1sL�

���=�:�L�h��T�2��5��$]L���+E�E�}�������	�d�c -Y��5IɣY�t�9�����F}6ޏd��o9VhG���R3y�hG��tp^���i�_�	����Hu��|���*��L���mժX	���A4�X�Pk�W�9z����5;��&8��J���~��er�aW>/�T:�����L\����?�������{Z��'�|�O��O����D�����:@�ӇJ
=����NK��B?�~����=y��M�T,��V��6j.���jul����o}�[�<��������������0�J��;
�~��]�[�y�2d��x�0f-C���j��R�.p��Kª�"���5�Z������촅J���Q�٥�C(��X�VgZ�d��~��ab��>`W`B
�1$�Tj���YP�i��n�0*-n�`#�%�mxa?.|�l�� �/�LK	$�V-��+�D�g!��t���"/7K�T��'�l�Dn;foa��~�pq䈷5�hw �L�RJӮ5�>��BI��尅D �6̲����du�݉�؟f�y�մ~}v8U�*)�����+�$c��^/�w��2�S�L(�0����TBL�i�:���-�:�4y�z�F�6���P�8�	T��U-�r�ӎ�>��[�94S������`R��ɋ��E�kC��J�H�u�줋�uY�6
�]������w8 ���9�3==��0��w��(�x	ݙ�Q<P@vr������[o����\�R�Ώ{t��q	F]����p��pQ !6l��p ��)�s\�`>�(U.=m~���T�d�N���Ν����d�ҏ��w�}7���f�,I �����e& .�{y��ٳ�%L�:P����9p�}�H�- �Ak~��h���;{�1�#~�i|��O�<�K�cǎᴘ1��>��Da�+�4��O,..���k?��O/]��b�tz�|'���G����~��<��C��c�Tc�<���ƾC�a.]�t�'�sL `����D�\�ʽ����`zj�M=����<W~F^E�hӰ���m>�3�h��?��^�Ž�<kN�$B��n4�O}��Ņ9�ЫW��'(>qZ*���~�L�M��߲$�����۠��k~v�����c$�U9*��k��I�.��t��_������5=�+J`��P���oI��L8)Mՙ� ԩ9~3kw!��U�f��LB���Ҋ�9��`��&Ӂ�<�J��=�3i��nn�;]H�j��4k�{�������j�i.����L���Pb�[�3�Q����	�ؚ��}����H�ۖn*˱G�x�;���qyެ7���j(l<�߸�?�����>���H�!VQ��S�~QTCw�����^*������3� :chz�(%iQ<��{P �������N���c��1pR���(I�B�jj:��^��u�ԕ�׀���s�U�pk��Z�ߜMX_��I��4a0�T�TN3���]d�� ���"���I���8�8�k�'&+Ss-#�a��|�����f�2aw��`l7�cj
�k|���w�(B7)�R���m���nGvJA�{�')�^X%�X�Z�U�U�"��t鱏?Tkkk�L�HY �[��Hp(�<���k�'Xg����$���C� v��)�U�1������DG̾�OL�P��q�I��4\'xkjL�������@H���ݑ�!���o�-���B�3\�khu��X�
}�ݐ���+]��0^��_*�[`Iz ������G�]��jB	��A��ށ=iI�J�$0j3�bGN�(p�Nv.��n]��оg�>hh"%��!�eP) ���ϝ|���֟�����WL˟�ɟ��������.�mNT}��O}��ÇMLL���� H2Z�Y[��?��?|�������[5$��녰��d���xcuUb&[��������zc2JM�J'��t��5.ZY�67��}��ycm��!��X�95�aM�n�n윝�n���U���;WW���+��Ò'��j$�D������(s��ϫ=�K����CC)Ѝ`*Ukmm�R�k��_��"�����	�<���o��̋�\J
9�~Ri4��&sc�V�X�����D�i��R�c8�\�5������k8�'��tcsm
�*��[��K��u�GP��2�)�8'���mw�''�PY��L��ҨT�j���Φj��H�deymjr^�h
�%̛�VG�v;J��fQo �EQcqaf������qc2�N��A�b���%,�[[���^4�R��dA_�pڋ��)��]���?����U�p�: V�%�l�"��LL��?��)y ·Ь,��{����~�=�]G��K/���H�T����y"�3���x� ̠�Yu��+L`7� >��*��7׮]ӕE�E�����>]k���N'����`7�7���k,�9	�p��  <�� `�҇�é0l@��ׯ��[�h�I @1B�?��	8����Z���F�b��C|K��Wǰ}����O
��  `��H�_�߿�O
�.:~�8NH�q�
��� A�x�"]k�<r�)��ԧ>�\�����~��3NB"�v����	f
>T��w�un��H��y���_�"I��  ~��^�u� ��E83`0�  Fzᄬ<�q����`5n���p!����f";ﱽ՞��Y]^��*�~��q�<��6�7֗Wj�VB��n5RE�ډ(�wΜ�p᬴8���,��:v�%��Y���uϋ�{���6����A�N��ܕ(�p$M�a��4�4����v�y��N�x>c�̖�6�<H:��Ĵ����V���5X���z�ۖtbl�<L�,U�r;�_N���! ST� S:Yw�@X�F�ඣ#B�2*%Ր>��ƵjЬ����եk��SӍŇ>����\Y[�v;�I�����D��=^קM+��DؖʊW��0L;� �瑠�/rP��@��~����<��G
�P	RS31ۋ���g/\�.�=��lS�A8B�=$��F􌆦�W�p�Zq�B��J%��B�Q	6��Q�w��6�V��Fڶ$Rk����߂��Tp/*2<2ۭ_���t�j%�h3�F���<1�o~�'��L5R4���լ'q��0^�>y��>�X����z���	iVG�"zv��6
{@�+�n:m��^Zզ��P��=�4U �K�$�r�ב�P�ecP�_��R��Q��Q��L�-�W�V˞��ؼV���kK�<x�4j-�V�97�+cs�����SNI#�����z��<E��]b�`�����Q#���V��4��׬��WN+�k�����Č��TR*�m���@��V���IH����vu?�f[���4���j��`ǃT�g���&�7�OaB�|�(�8TqUB)d�aK�B��]؍���ϔ�N��Ɔ�L��6ђ<�n����c�V�&���dHyy���\Q��16�6�׿����?�����Y�e���w��sϵ&�;w�>�>X�T���-+��^�1���������_��'OF����'��n�D��~ 8��Esx��	�Y_[�XY޵kas�}����v��h���~���Z��s�1�t�R:M4[E)u����W�.a]HMl�4�l�@�\��T�W�\��^�x�����8KUҢԧ���L�ν{��5�"�մ��j}���ma˒ŢMXn�J�]1�.����ɵ�7��y�k��Qؗ�1l����,r�"�E��{i�2����D��W
Z_�,���ݻlBFq�B���4�J
����-�2�<��n�3,ߴ�(�V�	t	��z��L3�bM��(51n[B���m�(��6��1CU����0�q������D͝��\-�@iІM�&l��f#P�m4�ٙ)�47YҨW!l-�\[Y�R.�,�j�^�K?�ͭ^/�h�&��lX���3g���M��%ALKK(�O�~��tq�e���������(�"���"�|lי��~���c�{~��0�tskc��TG7ca�4�s�%CTWڑIJB9�$�9� ���o��6V�nw@!��z~P��xJ'lP��pW=��4 `@�={�y�O�|��d:�8~��a�*��|'��I�i��4����HP%��[2�*���X��bx0�Vؖ
/��w�J|#��
_��書.� ���	l��͡C���j|��W����g�\��dY�Oj5F�06|�3��˗/��f4�
��s������ Z0�Y��a'6���,;z�(�6K� �fffp6\?g6Y���pi��|����~��MM` l��/|o^x����a5�<d�`�>d���y�\�?�aX	���� ��-�	L%fi2�Mw�R}�r��Tťɋ���՚�-4�+˫/^�1� �Q�����*�I:���Ӯ
AY�Qb��CN��9ݮ@ֻff�9u�ʍ�(�T��}�YR\/;]�WJ�pʶ(׊���Z�0���t ��(��2!�:����*�����j��In�sUr=���/+C�V���Z���i��eB('��J�b�@j����� ��S�oIJ�����Z�Rh*E3+����fP���}���/��te����FsD�h��fwV�g2q#�1�����6a-c�cح!�0u3Gl�a%�0���Iut[�a8Ȣ�kv���:�Z[_y��BU�Rn���@
�YGE�
3[����2e�������͛707��U�|��XY�5�Y��e�Or��i��Ô?s��#���L|����F�7�c��z۵�0l�X���=������������KN�
co "9xQb��B<�m���iB�#�!�nP�.�e�2�M�S�y��T* ��K�/�j��>��Z.Mn�תB�f���FiWw�'�5bsQ?�S�:���Eemm���{>P�<O��%��
Jqx��e��-�!K���d0COƳ+?dN��������0��)<�b��ư���3�e��=�-�瑤M����+jd7�D̡�ǳ˂�D>�q��q�E�nX�D	�v�{��������K��m�[gB��?�(��� �	W�Z:D�X����T��|�]�ʓ�!I�?ph�܎�0��o����ͳ0��8	݇7a����,��!u荛7�E�+)�4���믽����xj���'`V�S�'����̔�
;gmv��b���Pv������7���Ͽ��][��mk��Am��|	���*�'�p�e���Q.��T� ��k�3ѨUM�7��$��$!L,$�#k��Y�	�S���*�#��U���'F8�l,����,���,�i�|AU��{��PH����m I�� �S0Si�������6;�0��������4̈́�V*G9�:�yKMHS�D-�(���������/^x	#9v���������ƛo��li���{��EI�>&��=I��8Ry�i�d_�F"nm�Z�)��� ����l"�ť	�ⴴ�*f���"H��À��X�#<������i���u��>�O�)��vm˷;a[��㔢�G�Z�P�N��P;�ٜ��k�p��J=e����!XT�˛���Z�[x���f��� �A`������1_�z���ϟ^�Qa��aHs�_�Rf�[\������!��u��{=U�fm�ں�*���,	ǦGG0w�Q��*�V/ڄ��Pȳ��GS��
�A���	�( E��K���&�Ν;Y�?�����w��1.1,0M��
�5���V��1Y��a,;!�5ɲF`5?�`�a�a�I�I�c��7�@L�S�������!dv������?�9�	����|饗4̃���}V+1���r�>���������p�wr$df8�?�HJK{=z��C�g`B ki0�K�.�#'d�����y`� {��p>q!�jp<nw��⺸:��TC���(�Hc@66C�p�AƉ \ᰓ'O���Z�e1n��KKKD�.4@&�HLa��������s|�Ye階j��:���;�ûv���A���r�W�����²�Ӥ�S�8���hg��N�'H��X~`5j��V�^�QzɰדrI�̝,�*$3�~U�B��d)<�R����rǕ
T�ly`VU^��Ϩ�R���@�փ�����y��X�z=��J1�*K0�\����z�a^F��Qi�RI3�n��2]�Ϥ�Ep���n1F8MQ�y�Ir+jbY��,ia[�Խ��KW�^��|�}��*��T|W�JS��ZB��%�����Bu��6`$@���Х�(�������; ���N��p��N�^�"�oN4�A�(��L��ɢhT�p�9�b�]�A�˾��";8`�����3�af�8����$�	�R?*۷�(CY�+`\(ŝ�-(�]Ҩ��a��e�zo�vc��kqz~Wkkm��啺o>���wX�]8�{_���~��<�����j\�l��6Va24�%����R��aY�e3Ff�"Q��RQ�q09P�M����ͳ\EF�8K,勧e���n4�E�ન9K
�S�dpD[/J�,-�L����*�d�dI��I�ޅ��[�#�	�i#~d+�)�l��;|6��ᱠqhꚩ���Ǐ��/��
�:�;
a�B��O�U鷾c�H*��B��S�NA�}���e�_��Q��d9&,�sHH�mQ^QC\��F�a�ހ�5L҆$dІZ^7d��ӵ����qZ�qz�m=3��5��{X'�2l��YZ֪5׳w��4�*B��/`Ǝ�w�'v�{ʳ1l����LPĜ���,q�5KCyƯj|��o	b~"N%�?��π����z�)�1\w8���K��մHl�u�����~�w����[��$�잒V�o1.4��Ŋ�	�����Y������7M������cJ&yF�?�)�2��ڪ| �	+�V�b�d�ި�1&iبO��@�&�8J%~��39Q?~�6&}G�]��wO�R�L�~����uiݦ��jQG�&.�RCbALN��e*#�.���.W�/]Z�7n,K�DB�����?��㒆lJk��L�v�[_��	�k��uF-��>q�#o���鳧O�⥷O�9t���wݳ�����x�����˅3qƶ���ks#�<������E��=��|���S��ӧf�jo����f�H�r;��%v�	U���-�҉���b���6s@�(
��[�~�l���Z�)	K�&s�
��)�2�Z��
���5�4ߡ�k���=��`Y�xj��7����)���Acc�vk~箅���Z�ͭ���{�}�G�/���7�����V���-T���3����M���o�dyg���L���jW����@%�Qbv����p H;K�aH'�\��R�dÊF�9����ǻn�VEz3Ӎ���I�<3Xdq������wR Y�Ҡ��%��[���x�l9��!�"ï�|����V[��[�O`v�߿��&>~H�7�?v#et F3W�d�Y�!z��C��?���˗�B�k��LS��}����U�S�@DP����*��7��C5��/}�Kd�#G�r3�d)?`���0�ر�>��@0�&bcY�j��0ǌ�p�{� !t�{��{�wXP�]��Xc�]�����йs��o|�s��4��*��p���M~�	Y(pB�-�qB|x�=�`8ng��y��Bq#L[g���^�T��������D�9s��R�m+�� J�LQ�`f��\H��(V�K��p�smS�nK�W�6��/�C����Z��X�K����Rjvǎ�Bj'��,S5#��ԅ��"��FFh �a۫$g��޽{q� �ȍ ov�	��TQ�@�3���	;c������cMի[0�D2_X�%8�F�?�*��G�/a����`纩T�d�[�c��"��3� lL5��L���nŮ0L4'�(����$/�+�_�T�L�T�'s[��6��A����C_�T�0M�`�7l���m�B-��(���^�*CǶdF��RՒN��Վ������ "�%�
H�H]O�{&��Ыn������@�b���T��c��Ӵ�-���Pֽj��A�V��2#2�87 ��{�#0b<o�s��g�����k��"QlCWl��W�M_�n#H��`�$z�
׷��@� ?�ό|kk6�4�؆>+����Lj��9��o��W�c_�;��+�	S���:�
@�p�f����z:K�vbk@�E�����rw2ri�Zi��f�tK<�
�\�ʸb�K�mi�/�1~������^'{D�����젥��/��!���,6#d,�M@��������z�!�7i�h0�	��*�m?��8����v���6w�*o��k�ISx��th��@G���#���04������n�^���X!���>����ylfn���Z��{.�l(Y�ױ�v-�~����M��ͅ(�q-(��YIg6po�~
�W��
QJ�ۖ� �L~�-G��ҽ�^���o��xL���'>����d;�P[h��D��Ћ���_��߾��W�����*����̯�^T2ENG��4\�bfy�z�K��ի��7�}���D
�J*�#��j/D�3��� �j�:�v���j�V	�rӨFs�: ���C��[���<|����:��#w�߹��ܹ�VVWI[�]��CC\MO�+���y�QkM4`l��/�J�)�\�����_
���s��������뗦�v�Z�{��|�?��>��o}�;������~�ӟ������Yؽ�VD�V=�!�my�@��%�v9����j��E��z�s�BP��O����!鷋$��9�G����R��W+8����]����3�ACֽ���.�ܼ����nؒ��hV��%a4��Lz�a_)-qi@Q�þ-rY ����C���5!���T��=�e1ת����T+�8��k����]č���s7O����~���<:�B�F����:�m���5��#�p��<�C߉U��q��Uq���
����b���̜eV�:�ik�ll�Zu_���&B:}h�g�n �����XWVV`��2���v���8e��5B�*�����.d�S".V��0���n`�^!�c����x�P�Z�C�qI�NyAW�r��P�ϡ����ܕ���E6<e�Ly�&�}]�z��`o�'N�w�}��� ć�9� �����;!�q�ݻwCj }�_��g>����s�\:	*o
�ɞ<|Ό�AJq�
#����a:tH�`��I�6bN]��!�eH?�<p@rd�9��9��F6BT\�a̐�X���˜R`L�LU�|����_|�ͿIC�AB�aZXJ��n7����ַ��g��P��o���o�`|�3 ���:QX�RANMH�f��]G	�aӈ`�u�	joO�T ]���M�K%�M�9�}3/��bK��W.�Ѕi)},咒W �G�-�Xvw �%vy'�P�t�X֧�O��0o��əi��Э^Wq7S�~*����;a2�-]Y_YŃX[�I�i�Xq��R����P����'*�S�)�j��=f��Ͻ	����%9���Z�_J����R^���f�����N+umבt�4!W��lP:���\ߗ0�J@�eT۪��B㝠u�\ih�Y�=��6!�ɮ��=H�.��#_ُ`��֬�{�F]�IՃ@�L䆡���� ���{��e� ��� M�*ܤB@���X�F��aKd��(2�,���9I�Li��Y���f�X��Gxe�e�ٹ���[q7�y��W����m�[X-��4N���TUJ�j�� �5{q��8G�劂R�0�S�s66�X��X��i�ȷ��Y)[r>%g��Ŭ8m����J�"�T�tLU9T�a��4/h����(�,+Kŀ+��@�a¨ѬO4[�7V ��<[][��|��I����~2����~[���������Ly2�*�2U���uHrL�믿��_������m(����!���?��G}��ѣ���޽{�-~�%�A/���>�� ?�֏�MǙ	�B�4�䒁���jP2i'UNY=H�@�k�t��g&" �]��u�a�o<Q���:���+/����?�"�]j��'{��'q����K����>���W/���};1�o@}�}��=��̦VT����!��+W�ll�]�t�T��M˶���G�E��,�T�0�Ê�xQ���������.��d~��
����,x���+ �_��x�gO+�إw_���p�5J�G�B��s%� . ���?��{a��
<�e6[�?��Ζ4hN�`��m$I811�]#~@#o6�}���4����͆�ф�T�4��ߋ���&+䓪���9(e:7�P����7��Ѩ7N�����C�Aqm+yk�K�k�
c��TKy<+�4�a�1�5|���]CTk�dk��	��o+���c���cG^�W^y��?���~����z�O>u�FHJ2|/�vi4*�2p3φp�w{vgk��nIڋ���F���Y���^Ym�/���|������9� e0�Mw8��2�}�yj��n�[���N��+�����ۃ��U0UUA��O���ptn)/�R��Un���	L�0���I�OO.8phaa���ŋ�}㍷�]X�ꄙᗮ��,nG;�{+ؘ�r�E��v/R��A�I��' ��{n\��n'�z-.Ӫݔ�"�>⁓k��'1�����0RhtH��ڠ+��B��W$�Vg�fS�ט�.�K�(�>�<��:�	�����dq'�D;�xI'oS!��WR�E'My�DÊe��Y�H{N�(��e��� Ň؊^��(�#(���F�W0I̍�إ��Q?A�`��@|��NV8�7�|-���i{8Kb���WǏ�����p�	�(dǅ�[`$rOSmX�$_��WN�:���ӓǼ8]T���w�.1��웄O�ʭ�S9`���ũ#�����vp]��3g��Hj����^���d�ԝ;w_��ٳg��pQ�xFrX�EF���q�%8��Fx��̦���Џ?�D	b=�~qZ�,bK%�#�#�7~�����<��C�9�;�L2�-pQ�=0?�P]k�jE�{���D��N�y��j.^���F�	!lIC�܂-�f~ of�)c.v,r�J�c�n���^��r[�$,9={���VU�O�e�>�^U�"�	`.�E����MW�1�U���Gv�YT�Sݙ�����r��(�]If��J�ޜ8z����:u������}_��_�ܳ�Z�p�$���%�;��EJ�#��v �S%i)hr\���y��B�l`ɹ�@�kø*����H{�aի�~��ŃVkj�1��W^�ۿ��|�����?P�׬ٝ���+�k��p\�Eb���U�5x��ٸ#Kq��XSU������%���E�)�5,i��)�;�N%Z~�r�g����iq��V�fVn�۹���#|׮����������V2�HX�I�5�݂IAV`d��X�K��ԅ���(+����1���Na�K��)[��"Y솝�+�XP~P��(B����[�<s+����m� d����
�Y��CN0�*����.�g��m1|����H��,�25;5��`��(���f�1751����o������(�M�%�mM�,.b'��(��J}�������]R�)���<�Y�A��:>�ֆ�C���%�p𴤰N�i�+ԕ����X$�� �Da`$w�Lu�<�Q�@�x���"˶9�u�r�f�$�a�`�n'�"o6&�a67�l׆��P/�&�MM�F��ƍ�P�����T����|�;�<�4d��˗O�>qG���A0�������X���RSqP�ʤ�|�w�xC�@�#Q�ҫҫ��0��m�v���Z��i<U�ݍw� ��Պ^o��֎����j�|���_�O���ڐ���Xd�S�E�>������u8T�9����?y�'N���=��c{��U��|��~�/��'?�m23\�Ҧ��mV/�[�&a$�cQ�a�Y��|����'%m���аPvKK�U��IR�8M�!�`�7�B�C��D�YX��;��?���x�j i��L�a���k�c.������4eD� ��9�F;������_�v�?���+KKW�(���t��/��F�R�T���w/^�~ciǎ]����������ef;��F�(�`ڞ���R�(�<V����}� �_��MI�7-������O�9q�o�������<+u����P���0ɀ�S�"���Xm�DP�^� �|Fy������s/_�ڍ�v�I��[��o@Q��ְ���4he�*G�5���l^�P1a�J�0n�a�1ٷ�>����}�d����7��W����%5%��1�+*�_�@e���#�q��V��NO��v��$��:Y���U�lю�=�<NE�Дk���յ�ͭ,w����C�
��r�磗FA㌢��Gh%1 �U��d�I�7�?��,m^B#/"Ӕǔ�O�s�Wc����[��0��`B0u�!�E{�1R���	�Yp��8l`
��D8X8!LpN ۀ�uN�_�BĀ�}�]�_��0(�{�;v�~�:�;4�[o��qB����/��"�Ο??�^���t��t)���˲�WǥY>�A2����x\��v� ��F9	��0�s� Y����߬(#�% 5��y�
�7�3�x6��嶊���Kp�@���0����0qEh�'�#|B�B�G�~�@a�Й=��:ud��N���Z;�d���2��Tz�UB0�<���z�7�D��0�T��8��+��XdY5��F}n�UkMW�=�3b7U&ᶺmU,.FL%�B�S�7���G@�0:]U�F@AC�&��K�ҥ��?x�ͷn�X�\�PN���"W�^�ެY��I�ޜ��v�$��AK:S<[P���5M_����� ~ 	 !F"E膭r�=��b�'ss�Iׯ^{���[�s��{e
��حFszrҖDi���T�H��97��'>��l�e@��[��T���{[��I:����IA߿�2��m���f���ذ��^m��J�
�U�/� Zn*v8�W�M�ץ��KZ1*��|O��5��@���0L1.>ÖV���.��{S���@!�X��*nui�iH3*ˀ	V�����r�	i�fxs}%�W�V�%���+I��|K�%��9?��1�����0��t+��S$�XJ~�ByA�7�M�����RU��.�e;W�
̔.1dhX�TkCD6����M�M���^{���k�-�:� ���y�/|����-�	�33�b�@"��W-b)^�|f�����YiX�hA�|k��v/ޞ�9�N� �_I� �4<�"�@P�ٟ�$����,�[v�ͧ1'Y
FE�ntC�M��` ���hHT���<�qچm�����$���[��vB��"��Ӹ
�;t�����ر���t��*C�D�b�;�������,���1�Y�Z{��/d6:]#E�,�kJ�����q62IpH8�+��r�ԩ�;y�]w9r�՜�8����<� �(e+R�P�B���460?��!��8d�ٳg/^��y}u���Dq4����{�ηC��Vg!>_�&�#V&���4c���|%#�f�{A���-��69mp!��XoOLM������?�{����D��y�����233u��QXg�
���*��g'�f��<_|^3�3��F�*Z�b3n1�����v��01�7o�u��ɓ�߽ ���)��Ǽf�w<�8�{j;}�.�K�E���ʐH��q�]\����	$ba߸qac��ю�"�c���M��G�7�B�ާý7
�Lo�c�Ui��c�%t�F9*�[��ཕ�<\���F�?[J��2�{]�'	)��:�@hB�m
��f��Z�#�ޅ�n��4�rZ��|�dR��W�L�,L�(��V:�xy"#єh�`*_E	&3��������7Aהx��V�tX1��V�}`:�l�5/ǶӚFG�4�&�*c�̏'�y߂���9-DtJ��21;�n�=�F��`��h�/)�H�͎�a�о-�2�L_ZZ�5�G��Q�sv�<s�q*6��ia�b-rg�|����P���'0�g`��8 bb�6�	�X�X�i�|�Ն�bxW�^���{!b�O\��T.F�Sڋ�A �MfP+@������ϔ�//|��wc1H��tۜX\�y�쥋)}����%��s* ��3���b�FH.
�IZZl��檥�JXB.l�;��o���@Bm�*5Z�����X�F��#��X�vБ8	Kht���\#�a֨�K�y�ڰXC+
Wa!�1�ҍHe��v?10	n�Q���ۉ���E*��Z��a��4Qd�2����Z�q�����^��k++0�����Eկu�A-�h��Tka���ݻ�8t��+2�v�'Hsjڰ
ϯ�A͑ƭ��Fgk�0�\S� G@�������%YR��'%�*ըU\����	Z-��Z�ދ�L�����._�y�!�{��]Xo�O����U�O�+]���"�"o�ǎc��� �}�i��E�{�)��Θ��F�vZ��ǧ�F���`�\:�C1�J 0)�bT������W�r��
�eK�qx���r�0��NRgPS�L��-��Dr�$�UJ�Fb����6`;�gNP��[��ffY��cDD���ɨ��YU�ny��-���W���s�� t�ɱi��0�	�ް�(�~ 8�:�*n\������� ��T5s�}z�x�T{.a��ߝf���;��ڽA�۵67Mũ�h�0���(�]٧6{J`YZ���ǜ.�$�i�sTZ�+P��[�b[2��_�Ie�HU[�dwTM���� ��6D��c��d�4F;;;+����f�$f�{��HSƀ�g6�fёvѡ3��t�GUkU>�m�q^�mw7��FW�&�c�=`����mGiw�F;-���v���I��Go���ׯ\��������Z^������V����:��= �1L���׀r�x|��''�IA�s����o������Ϥ&��4!ZP�\�9�/8';i�+6��}*��b����b~��m��a��������� �lD���4>Me)��2���N$b����B���G��֌�+ށ��VVo����f����0o����9����w�]������iY�&���3���W)-�T7��U�k��»�+<Qg�p�"���ץ]���*>��o�5,���V��5e>;+y����,7�Œbы�$!�QĬ��+�["+R_t+|R܂C�3��C��ݰ-)��2�*G�4�e�	�q�@�:�OQ�΋<3�c㴭��E�	ŏc��bJ���0��\):[z�:ٯb5ދ���-n�Jd��
��6Va�^�����{�6B��8�0T�o;tS!��r�F�.٩����)k�(񀘃�T�\��"�Q&�;��3`���r���#kYv�_�4�k"�j�۶���P�yF��m͈���x+���h~8��m�ՀeB�+%g��ʳ.�Y,��6#];-*rX�w*>!�"]5�R�afH����h5:)�p�/}�KO'O��v����ÅH�0�^ ��Ç�� G��9�P/`�Mt�#'.����Eq�9i�o��l�t�w��a`�>�9"�,�}�^� ��^i���Νc �C�>��1Ӓq3���A!�
'�;~���˗1$��uq\Q��C��vp]����&�c��6>���>���>��Ɇĕ���W�m� U�)���1<�ȥ����t72�
8���8���l���_I�h�O���~��rtѼ��f����� Q�#���cĴ�}{����D�*&�\˯W���Φ�Ep�a6@cIG9�Q$��}I�w������ڮ}{}��X��;�*�Z�'������7Vv�i�[��n�(_�I�^`W��*�]��[���J%�߫�U�E�^{���]X��ۍ������CG���e��Gz}uM"�FIW1>�*�y��^� ss#���V�O;����� �p`�Ì�,/<��I�"�b����ϣ9W���+��6/�E$����1$��үY
���Ö�T1����,��@��?d�{{B	w.}R���y��O��� 8�i��CqV�LqAz�v��k�asr"J��Z���Y�R����˗�x�	�2B���*�<�6և�[�NmXC����_	Tђ,]ۖ�U饡� nk������@�$9n��v�� �Xg���pD������'iT���{��G]��8N[�=;�1������x�߉�eկ�TZe��F[�&V�#N���x�`����!�۵�n����kƻ�[W/��`���6�*�+6��XA�v�ǅ�2�"b'�Ȣ�#.�gp�W��{��{;��x�*�!KU��J�R��vt�Pc!�����M�144��ō#1�%U�+d����g>�����;��fgЋU�^���=EO�0f��&���z׳gϾ��ۺ_n0�=׻:~P4�:M���|���o/^��ŧ�y&���(�ęٓe�BA�+=�
U���L��~��߆iqp���7-��4�&���0�a/��f�T?:O�,N���9����=K�֪��<Մ�TO6O����>����A���B���*���v��c*�n��9�=G�5 /؛�v����W�n}���t��SgN�z��������!���Q����%�Ԓ(��]mT&�-�$��v�rm}�V��a�*��H��Ŗ�6��"_ڟ:Cns�s��Ͼݪ����9d���z��s��K�:�BC8>��[��a.�����w��+W�����-;�3����7���Fh��@�I�H�"%R�������F�*�fʞ�_��*��U~q��e?�d�дF�(�,H� �� t���{������9��}n��fX�Ev]�{�>;��Z�[���ܳN%�X�@ ��q'k �9��o�<�J��$�b�;�Be�?�8���_[A�B#%+��MŌ�c�q%��,�,K,a�A�?:qǓ���̴Z>W��<�+��ʹ�C&���ˡƩ@��CS��ҪrΕ�����%7��'��.Y�s�rN�J3%��DV�m�.�%6�ܹs��v�6�	�.�UH��!v�c����	N�����᧙���j����� ֓;�8"�����C={����sw  K1
§?~o�g�ܹÝ~�,s�rG_��� ��M.��->���w1s ���u�8��,�ģ���$�u�۲���:�L>���܇�s����`�!�.�	$/�\0�r���k���q>����?��O����w�R�U�_�,#Q�w����9u͋
g�*�̑�Ҩ���!�_�����G���\֊�J��L	ᡷfg���O�v�#<*܈�r�e�6�s,�<�M�⃙ȵА�U"ćm�����(X��ɕE�Ȃ,�{iJ2��VaY31h~�!!�0&rm��/�/T��x��#㴅�}r��G�f�-�7_���."I�k�0�a�t�IS�����f÷4�	�6"_���m�҃8�����,3j��	�F�2Q�:���l�ڇ��t����_��{���F��X���Q�b�9��E���>�ƳgX긁8=�u&m�$65Uf�?g�cCy�f������!䢕bLK�h��
.<V�1�b �u�r@"��ĘcY�\4�M��\L"�NE9q&�e�x�e���I��[L�I��5�ƴ:+O��<�B�I��a�|Mi���g����q����lgΩۋ3m��hx��Z�t���Nͱ�������{�O���;H��;3���ʉde�Q��5A\�����N���NLO�&h���W�)��AO�HT12�AŠƺR�K�)� �#m�B.�D�۞�#�.���}�cni!o޼�3���s*3j�Q-�Hwްl�7�+�m%o�R����hN��Ū�;�T��"9wz�D�D�w"	��z�iX�����>�_��Ôq�>[�C�P��¬��:`�T��_x���'%C#!y���-m��Ã.U�(���"�:�	�v�b�&;2Νq�Tc�)Hn*��Y?�,s�/�޶:s�;Z�M񳽽?�Ņ�43�� ��駞:}��ٙ���U���c��υCXo��~��Y`Q�
S�
{�s8�݉� �Sb��Q��(�D�.8<�����f
�07�<y���QN�1�eAI�iP��4���-�~�`�Z�氇w1�����o�����o8B��@�y"�e9�8�ScBpzd�8�������g>����������%���C��7d8�_�Y�Eg���o��������?F$���(���� ��KL�IA"�Tץ�3M�� ��_�l[.�������^�x�O=����Qˏ�������h�i΄�T��`�O�$�@S<�0��-�Y�ꎂ~�P�TL��1s��(xS�P�rB):���$�[�J\r%3������:��$:�x�R�ڕf��P�鐉
�����Tqׅ`�.TZ�#'l5,'����R|�b�$��*KCi|���c2���7�1��o�A����Q��b('^��`�� ��n!�J��0�vgg˲k��Q���F�F{��MF�P���K�3�Z�(��U�SiR���y��O�L�fd�4�UVY��:���l�%c�˶L��������vb;D\�`��Ex�J�Dׯ_�8r�̫!&`ve��eQ��80�|�̓�h���y�'�C�0
�Fܰ�����E�����   �� x���{�9D��X�o;{�,pN�}6=p��88^<}�4�2���W��k��� ��5��᯸R\ ^d	Z��C*΢����~a��}�k�����s ҰX-��� \��&=|`_̓7�j����')}�s�ÛQ� \�1�N���x��n)��c��X/�US���*7J1��L�3k�K���� f^�5�D��S�iwh%�Ao���"3���9� �1��RΤR;��T��#�\�G4b��P"�QJn�S���Q�_bu.�4�(M�,��@���<L⒒���23K-�	L�d�<}���y�Z�V����8��|�m˩�c�:.[^��<��z�,yڪ7�4���j�|1�X昞n���x��ǎ��6�y0��(}�k��?��ϯ�UM�g��|�o�,�nPo{�h�:s�Ie[��cl����D���˂x��H� L�L�wm~�����Ä{���Y����m9��Lj�0����]���*�@lmv bF���MZ�K��G�'�WL�� ��lP)>IhY)�rL�4���Ki��!��G|��^���񐇸�O~⁯���O�<>7������˯6j�c'j3��>����G�^����=��<�������҉cZn�g��;���:��+��B1K�w�� |Y�նj��>B��q��o0\��Ѳ�$������h�Kض,``[��܍$d�ub;,�V����@�v����g?
+��ͺm��%���q�!��/b�r���>��lǛ����I��J.�^e�GfЪ��S�ܼ�8����pD�!F�"�3�ȇ�cLrͭ4���.����#�reC��իܟ�y4���ճ�Cz�F_�s���X���	[�D*�-6S&Ȇs9�+b����[%K��$OO���:�3;[�XH�p�B�|W._�r�򱣫��<�8��h��|*�*���D�9�A��/\�X�#'Q��`p֏�h�h!��il�����I���v�ps�ٹe7�#��*���8N�&>��'������[o^���cȟVk��2�EY�ԅ,�XJ	5U�s�2�D	;eJ�@D��YzY�+��r�»;�)�L�#(���b��������8Fe/���������|��ɓX&GV�h�}C��\Vu8t��P�ZF��;���#����mн��[�g{��vtU��Ѱ[�sU��
�ƚ���������f8�y�М�o'T+���I|:�5짛�i86��Xx�ndp����ʽ��b�B@��R�Hy�0�-Є�.g%��mzA�"�h1!ĩ7M$��: d��n--�����'%"�1��E5u���?��G"��O�`�%A3�S��j�L���i�������ڔ���R�M�!���%�\��t"���O*��~q5�O(�S:��VNUidW}u�q$�}J<^"I�l�I�l+�fJ�"����?F�n�R�vK՞�j�S��)�
����766 Z`Ȯ\�c�_���:S���x^gJ%�$�g�N�A?�<��87Ƒ�9Ȥm8��a����.����ae&S ���c!n�����#�g��`�
 J���E�㯈���/p������`ނiv�q�e|���2y�	_�?�.��|@dEN�w��'�j�p��J);�K�\��-�~&.�?x���Ge�7���?����G?�9c����pB8�/���;z�(��1�&A�ѹV�S��	��|h\v��<�N�ɐ�\�J1 �:���` ��J�
��)A�C\@% �nW��2ga�ĵ�?�n��g��혚�$�l�z�yY�"�ZE�d���#gP�ZGwV�
��z�_
	j��t�3�`���I�֛M�Wu��>��Q����{�������-�/�����~�w�� �5���Z��7kuA�M�bn͵lc &��P� >~����u���
Nlcw�D�e��?�oVW�|��gw��~��}ay�̒� x V#��Q��oMP��8˲@`��ߩ%"��7[�t2�\bq��S28�aNF�I�U�&��	fx����wˉ��#��0�xg!�ZD*���]�Ew6�w[\18��D.U��*�bӥ(V� ��������
-�QmZf�Q\E�,6��?������!�!X3��+�Q@���bB�Y������O|G!�CEԯ�B��_��׼F����?��|9GuҪK;�Z��b�Xm�\��X5��Bx��\�c%�0*�#�I�)�,�hF]�K5��#4I�[��tZu�6%���o|��|O��'�|�ȑ#~���Y���[o������O�ڤ"�Rs;��̙4lg���Ќ����Rղ]�Ӫf	���ǲ�K"�í���t�0!��<r㢙mܺB�*�%��ey�Al�G֘cFҸ����~�-Re*i�,�L��S=r�d-������s.}K*9����r�*�dY�2�+�	�T~`�*�Br��N.c~?��4Q\���b#�6l���Iv���;�7��]�5����	 �|X�� ��
z��	-���'K5�`?�E�NU�$���+�7�W��çpv�o��sU7i�Y�/�����|�����~��O=�����,�J<���9(H. 9��	i:�%���i,6Q�Q�m�3p-��Vr4���/�Y-�2�3��J
��SZ�d�A0N������v���O�3gΜ9u�T��z�`��ܴ�	�X�ؓF�& <	P���;�/_|�����׾�k���/~}�7�~��o��w.�w��IY����$����#hW3�P|�O���ߥ�Y
~�"M�2u,3��?�/Q�2��O�
.9��t��U�t�	1�(����	^�)�Й���i��O��eB�<c:m||�2$����LCK)�+�5�a	,B��DaP��\�/��[j@�k�i��_M���GaJ�|�n�V���7ڶ��3�-�M2bjM��Z°D�}�A�!V�yAJm{9'�9���m�)��Lǩ���a���ɻ���*M\upH&r�&J��*i�v�xl�Z�?`�Ӧ�¥�J�UG�d��Z���&p,�D%��g�`ü��K����� � �����'.Y0�6���x'M�{�=V���e����"|������h\����?�W^y�[�pOΟ?�C�p�/_����=D���,.�:L���c2�5k"�N�<�%#��k׮�!8�g�3��� L*}���6[�U���|��L�)|��ﾋۅ��S���w��2B��c�%~��"rV�ß�Ύf��+����� !����W_�t:�X̔� ��p�����p��x��׿��oq�'!Bb!~:@D�O��b����~��M��(���!%���߫�$��w�9�F�� ���1ni�X�Ћٿ�w�p���jQw��������p@��eK!F_����}JpƑlE���a�����1�,/!�誐0��j�)�X�E��E	eL�0iԍ,�Ks�O(K0�o�����{燽�n\�������W~�W~�X���_���k;%h�rpsa7���8k�̎��GW�f��������\[�wl��)�����|��ο����No�w��COZ�VӅ#�X][[\^�b�qZ���c)w˂1�fHFA,ۅe�8?���"a3��YF�!1@��o-'ь����S�$+0�]u�j
�T`&hc��	�h�Ω�A$��:$�����b��/`�oFQL
d%@�����Y"��Т:g榧ys��*G8��-�]���MT�X��
VW'M�4R�$�5l�$�(ö}�QX
�,�mΘLe��jd$�b�P�.���-z���B��~V6"kl�ÒՓM�A^�o�w����n2$�\� \֏]}��ǰ�)�7M����E/���=v�ѥ���^
^}�幹�p[�̴�HK�"�5h��=x��R4!�Ņ-/�L r��J< �^�C�2	rx C>bN��MJ�)��NX�L��rtV�0q�'h�q��A>;nf�������k����K���@vLT�5����$�*_�칐�ޕ��@�R��x�K��ɏWC�ː}VU�nw�����x=	�[� �$�.��9%>�w�2AYn���g@���awv�CP'�[܁��Z,��#��n�C�1���ja��K�`0H�n�|�l�R��?x����O/-iw�5���޺u����)�%��Q�esa���)��P��Kb�,s����"���d��)2����;5tŲ)A&�5I����{� $����rL�����}���{��Z=՚��:�1��̻�p�ݽ� ���_����o��H�O�Z^l��đ���͚��ׅ��[�T�����G����b���y��hv�E����¾kZI8�����^(���2+S�B�NS|�	au.��puLo��b�+Ih��ShZ)+���@4�\��JZ��" )��1�P����_L�$��	���$%���rt�����Z)
�:� �Z�|��[]!Z���U��5�����`�z�%IGϣ<�Lʋ�H$+W_ɺ���h�;��^Vqb�ô|x�Hd��(%e>�DT�F� �Z��<�Aڅ��驝�n��%@7�A`�5 W�1�sY���j/�/��Qx;��p9��-v,S�F�J-ʦ�J�2K�^�qY��A�L�U�%Ⓓ��qdg3G�2l���rTTzh~�KLm���l�"we�j��$�s��P�p��K�8�;�^\����<˘A1~�����u܁�	\�`�!R�m4����w9��a�/��V�×�X�_��c�<��zv̎���|Jܮ�
�8��I83�%��7�|��.$�(?�g�yF:��c���8��^{��p/>�u3����7o�#����p5�'��)�1qn'����?�3���ĕ.�g<|Ŋ�a�jBx�c�@�81\&@��_~��w���G`=q	x(�Tx΄���s�����q���d��yM��4���n�Z�l6LCx��u��RGZhe/����%E�[qͲ;s�������~�[s�ۼ���`f~naq.ɕ���ѓG�����g��8�ߍ�#<�F�tۖc�`.�a���l��..^���s+�IP(E���TD���!5m����qZ�%����×��ȳ����m���
 �mZ�{��w.\��a��oڑ^�q���0���m�N�=� uؕ*�LW��STk6`l�ǆ�Ԑ��Ӵ�lw]7d=����ہA���'���ѳw����o��y�bx"W.\��׿�G�aQ�j�2㈔"a]�q۽��*��m�?P)�m�<eGf0��8�
��8I�	#0�Q��y�7�c=�(���E�4�p�h<"�P��v	Ӕ�8�!��B�T�K	�1�^�u���5MOD7s>�o��a����'�M7:�$M�|�&�Eo�`?S���'r�����;z�O�L�7�r�֝;��s~���֎��v��T�o���.��,,�,�s���8��ob�Ô�� �XT�q �BQR���)��5��j;�w<��얛����D�fQ�Y�����8%.�VMJ�����2Ia?5}޻��o�<��Ϝ9st����m�2�z�J�!���^���#g�=�p�����y�W�x�ܹs?|����h���P�,'0�h˱�4LF� a3EaX���4s�f��4jT)&J�b�I��d�PeܑX���[��q>��8��L54�s\�!�B�]ϯC,���9oC��Vl�̋�"�y.q�1��1���`��S+����!
�@�2�(;��mA&+��|[����d�ŋX!$!5<��ɕA=V��C1ZcnS�ۍ�K��C�qCw���Q?��s� a��|�6���[Q�L\�8��[�8��_[\�����F�	�6����0��q��
�<g^�������9��理�n�q�¡����<VB!lF>��Ӛ�*����������뿼uS���~tO�T�PO��$
R��*tJq~7�0��=/�48��U���C-�\_�FDף��\NYZ�U#`$�T�<EQ(|A�>��/���#$D�h�sd��С��nwo}����m]��T����~nqa�hQF��5�Wg�Z�{���*Y���d�/��xq��KR�.k�S�iE��{�������ǜ(�5�1�����X1l��q���M����tEf
�B�%�H��6U��!�/�1k� [Ģ�C}�c�G*p$�a�	����U'�7E�?HC�&~6�����%��(�4�Ώ��{�k7ǩ>��M`D�ĵl]�SSpSajE�/QLK�J��w����L7������(��U����;Mg�΍A��Na8��:�� ;v+���Hg��>�����kA)�p΃�A8�pbQ#�E`�ܱ�x���(g�Z�U�9�X���h��3U;�j������%��\C�K��ES	�V;��m~2ow�L( 	�Of��j�� ��0���N���q���:��8��;��g�`���/�N��� ���NXK��%��erq������\�_
s���������L�q�С�%i��G�;�f�Y���� ���d��g�>��#�H����_�	�������s�C�<��P��h�x�:�gf���-��Þ���ﾋ�_a�?�Wƴ�f����c�!�R�i`:Ʉ@u�7x�}��	����n�K%��x�R�CO���2����c��$9��v�"	%�]X�
,�7쏂a���o���Qda��$�x�ݗ^z�T��g�u��m[hFA?���Y�^��~���Q��^
V��q� �4*�	�e;�FA�������,��]=�inׅ������?�裸�^~�2��c��f8��L� ������=VþĽ:bа\�x��?�9���Ϭ̯=�̏.��>��L�Q*�}�W������0?��6Whq�k��'/x��_xQ��~��^���X[^��c	1�� �h�w��|iy�1���j�(&6�)����GR��%�H���d؄���\ђI�	�K.��F)B���xR��Ga\Nԇh�e�&���ְ>����v������b�?����닫�`��_��?����X��_|���ٿ�t���͍v���cgO�:����ko|�[�G����:~�8�<r�G2�����s�X`��7��]���������_��Y������[on\9od��Ң"bS�A���1��C���v��^�������sd�>D�@x�!F�=@���>��U���-\�x��o 	�s�[^^���X�tD��`�.��W^y��ɓ<�w�����H�_�a!H&�fr����{�^T�z�80�9P�:��{ݝ��F(��S��a����N��m0w\�f���|��_�ȕS{<�͛B�Lʚ�̎K+'=;��-�|k����:���H�HJʞs^�,2ΞNMI7���fV�D�c�|���V��u�T��tEI�^sk��y�
��'�$x�C����'s{�Ŋ��{6��3Z���F�3,�R�Kc℩vA�ن��-l�	��j�d�[���X���f��";�O�'�G�"g�3`r��f��5�''U�05߳�K䋇��pcs���B�>���p�۱}�Ed�f��8Gy��_���vaG��(A���i��Z-�8��59e(�/�I���� �v�s��_��§?j���ff�ka��q�S�7�o��01iݨ��ٚ[����8�(����Ͻ�����H�53u�ĵ�D4�4�xӎp?3ŀE7�tcf�Q��@���8"���=ķ�0�J��0� Rm6�l� ��p��n�&ްh�v�� �7�9ُu�j����H�!�߱��������5a�:�Y��_{���V�S�$^��c3�5r�����u,g��͗���[�mRM�0��k����ɵ��=Ώ2�$�-�)D�{>�f6�S�2�P��Vث����fG8��^EG���*�����DM��f� W�fc.Ȼ��ҖD7�og��ѿ�s�5�`�$�~�%,����̨�.�����䤝�cw��q�����a�W&ז�ε��,�0�L0ӚT��묫 ��.� �<�$����	ֹo�v2&��F�^ZE�gȖ	N���<��C	��-b fe���9�eAΉr}��^����=��b �F�����y)��l%�t���gYW
ny!#ZJ�wZ8�`��x1TYbىrI�HQJ
�/Ј������m��y�MO/���(�Qw{&��y�j�v���H�Z[5��2�7,�(�4Qf:� c�����n�)g�>���sϽf�i����u�t}��wQ�Va�ko��,�w�����y��{�fx�ȑ��93��q��|W�ۻ��!���	+K�Q���G�I��ȾA��;����X8t#�_��v�gΜ�����歭ް�*+GnݺAmʆiЬ<3����9�ő�.��ggg�p�S�L[��c>�,��J��)�4�.��j�P���e�LJ�P_T1S�)�,0�\�1��1_`�_�۲�Fi"q�v�R'�rfH<x�nl���(����/�w��k������^�����U���[�����;%͕�o����}��bx]8�/���'�_n߾����6V�%�������{[�����������P�Vj����K?'H���߄B�aB��f{��;v�|ὧ����?�̱��ť�G9��/~	�ysw[7ip����F��~�ӧ���qb88 =�L������1�n+�Ҳ-��?��?�����#X37n�z��W�XQ�����KI�'�-�̙B ���3���R�a�M� f��Kv4�?X�ܬNfٯ�����˗/s��r�� �
�v����~��� ���)g{d�k��[�eͩ1I獽 ���"��R
�Z=�*�V3:�'�cZ(��4�E�����8[����n�gHV;gٻ8�<Gv� �5ܰY��߿���2tA�Ǎ��0e�3�+�f*���6��U�QE*�D���P��A���U ����wό��L�Ga��^��ױ�4\�:��:�P������ao�0z�{��Cbu?�aZ3�0�*{gF���ťK�����|�Xф����2Y^P�^�	ќ����N�D2�O�諻G��4j���q��H{p� �$�����w�(�juX�V��f�B#�9�ɛô�à���t�o��b&�0�l�U�P�`���H"M
޽��y7aT\������JQy1Ӯ����.PY���u-o�U��`��d�D�k{��" 9�Ԛ�V��Î�Nd�ñi鞋~$�0�כ��t�᪶��j���v�0����2��p4�>r�b8ݴ���3��n�Yp��L�4gI����
AQHrX�(��(�Ƭ�<[B��c�v3�Ƅ��JUb�yK� Yb�N:V*���L�f�O�$	Xu�RF���8����UUf�*+�[@vKp��"�床l��$0�V�k>30�<�nV/���)�7���`#�8D����D����Ӧ�t�͏3pU�HSr(/I�`O1o,)��}}UɞOj)T%�%��O��	��G}�1������|��'����i����B��z2�J���7Kfv�O��d)!Ώrc��?�˕�&�Ǌ%�U��9?;���"��=;��#7�����&���[��+��p�Y�Wך��z�2�$�I�i&^���R��^l�I�,��yƽp�(�_\����iJ��N�޾�yg}����?r�ؠ>��s���dvv���D��좙�4.4�%LYCUT�|f�nH����������-�U���^���\U>���3rK5_�|�ʵ2��u���������K����X̲4Dz�+�0<�͉�C؛0��p���P�F1������m/J�;��T12�����qNK˜1y�I��D<DĲܙɈ߂G��ă8~l�b��.y�%%&v�V����gǤ��ʰ�S� ��6]�.�i|u@��iAp���(�!�:ĨО�ǃ���i�d���/�8�cD��pŌ[
��L�c�GV��n7Y��)��ۭVQ{��/��8^���ܺ͢�8�C=��"'#��ej���q�X?e��4
�3�u{Q�cXN��b������&a��xʰ0��\�%�-t3m���8��:�կ|~c����I��Jg���Y��qA��h�����S�"k����.1�*�(dK%��.\�njAL�^��ťB �K��pa�Ƴy�Z��49;*W~|�xx�N��>�P�8<s��/~�WV�h)RM ��ظz�"�Ϋ=5�K�hnܹ���5|f��;WV�aH�E/��2�>=Y���p�1G�b�Ѯ�+�l��+q���
=��R���>�d�k�E�Μ���h�L�6�\�t�)���������n~��k�TTi�ZG��E�#DlIQ�s �H�3Y�ئa�n4�i�@�Hw�-��n)�����zɤ�2�1)�l�J�p���mո�:�U��~Z���>���X����K��	A�wl�m[F�X5Yu�p������\�ǲ����&��<kR.��B7��Z��#F����M�$d&)0OB������d9&�^FA���X'�Ba"8(p����:�ہ��,�Јg�P�<F��QG�	d��!2]HJ-���LB�MO�R�q�*s���s0)�F��՛5��Ջ<���lhQҋR�Y��5�-�,N��2=Ӝ$7�WC��	���N`ȕ�
$%I��0�mg>�4�R���tt1��*|�-k;���T��������V^��'qf�q�'u
Vu\���w�kri��^�z��#K��k�*%~4�?
����d%]6�UM�"M^���ZI�6�U鳧(b�<u��	6�W�����$��,f��N��$��LxpRM��C�s�A�M��+7r紜ԯ^ �w��WH�Q٥��:_���)1��_��alS%We$�?��悪|?6u��R	)0
��ς��K�0�*���!��~�o���g?���t�ʕ��~��͛�O<�w�[����D��Y6Q�W��{��_5c$y�rh�v�g��f�ΏFf��*�x3�V��K���cȊ'�2)�����e�� F�7���3_���ug��������b�=�j�Y� V�v��m۩)��u�ǩ���o+Z���#yi<��s�nm\� ��--�ܼ���f�;��n��m8��}%)q�*G�R��],^�Pj&�{�酧E�������z�ٖY!`/q������kN3��iz�X#
G������۸a�*JQj�����d�3i� 7���ఎ����%a�w���i�te��\8��{27�g���*�/7���R�Ew�������3 ������ӧ?��C�N��X�t�4��{�\�%TjZ��ܝٕ��S�pZ��*vL����mUM����0��峌�D ��+;�x���u`Z�j�kcaP��T�����f��'N=���߈}���|��%�,)�A"��>t֬�c���;'O�<z���I�M���V�������;�v�h��ey*qg'�w��XE�����B2_�F��Od�Aܨ9u���]Z�o����Fݳ�O��R�H��~��{��<�+5,�E��{��b{k�+!����1lVDM�0�X]i)Gh�li���'RTc2��-�W�M�f��_l��R8�\���x�<}��F{f�{[�ܚ��FI�l[g֙���\��꽨�k�ޓytp�v������u��?��H���e�����I�3�s�n�8��TZ{i�eB�p��z��5��{��+�8�(��|t��}'�p���FIQN2��|���'�)�Vg(�1��k�WVV %@ڿV�YY]���% �y��~��? ����Ь�BOmv����ŏ�]s5D�g]�G0H���ƙt9��{�q������>wO�{8e�2��>� �f��i��5ѦA6&�Fܺ�O3Nhƌ;KM�j�H>Fw������c�N�2/���ג��cSS=`�DvJ�P�%p�4m�sM�UP��gi8,l��--J�a�6}xU{)i�c��U�Dk��;��������l��+��BOq@�T�E��S��>��'q����멣f���E
xШ���.���F��Xef���J`jF�шr&�,�Rհ����EF�o�(,ۤ˛��kI#�X��31�Ȣx�.ľL�P�;�<u+V�0.t���p�Ru�]��j��%{e��y�F�+qZ�ڄN�pe�&a���[ot�W�w6Ԝ�+��y�Q$̲��*����j���N�3��'!�ʹ$g�i�Zة��q������27&�֤	�JT{L%5B5%0��1��R�3��j�ۯ��TQ�����fXX����'��Rw��6��QL��T�L�)��I�nC�g��΍gr�G�QpoRU^��:X��3È�7iJ8����]�)ٟ�ũ�֐�:R�Y6��OUe�4ך�~r��uDW��T���pE0�ReU>)�t8�)�����*^�m�c���Y�^ÌQ�H�ϋ?>f��KC�1I %�xb���=!/(�q���P:H9)5L8�i�����G��>~j��wn��~\ZY}��s��Gq�u���n���߾q���T �J��V�^��.P������Rt����ǎ=�𩝭]��>T��H�Y��d�6l�������KM������U�̎�8�������s�.���/��v�ܹN�(�+^�v�՗^�sg���<���go�:|�lt����,Y�� �2@,�{x��ǉ�=��,	i����jmm�H�ӆ{w�:��v6�LEB�	1��Y܉����̀����ɱV�k��c[��&Z�I�G%J?��ZV��F�8����d�8�S�R`-��H��(��8uC�jm$p4�0����t�a��\�U[s��{2���x���EzA��H<�(�|{g�':rd�5���L�҅@񮫥�Ht�l6[<Ζ'y��M�*U���kD �F��b��ZYk��'�pf9$-�zD	T&�c�yJ,�������9�z����25�{-���L�K� [
�Q��f�ӃQ���l����F�v����T���Ʃ��0�E�VՁ"E�(����1F��"&��� ����;��/0�̷ B�`%�Y�={g������w��s�Dw��r�(B�\��؋/�$Cga�&�F��^{�7�`�3|���p��W_�ըo�ԩSx..\�K�G�f��ܪ`C�X��p'�VI��f��Q�R�YO��ˉ;N�qi�}�*��d�A��" (ӣ2S��+�^w�ڵk��=ߚ�`��f��*��(�Ƈה,�ϷLVN����#�<�g`�4˔�x�Q�o�����0\�ڡJ�}��+�Sd�&c����e�������!�>���$������T��c���^ 4]�Y���j!&$�	�oLa��!�Ln�B���BR<�3¦�6�\զt&��Gu�ψ�BEo<6c��0n��ߟ�&�K*����)�LZah45��:���1��:�c�ؚ䤇A`�<N���dI�䆣!���Q�h�_W
�nAA�A��^��Xe�h���(C��WLK7�F��R���j6�r�Ժ�CyI�m�?��lj��iÑ0�5�)D�նHȱ�P]S2�	�pk��90D��4��`Ԛ5E���h JQ�� ��DqG�9|�
��:5;xd�LW���;����YX��0���XIKS���҈����(I
t��BtC�G�q''�}W8:�TS���:g)��9j,�1ዬ�>�j���TWyU�j7�����SB������R[���Ρʯ/�Ыw��J,��@ˆ��l)�y�dA��X��dQB6�Te¹3g��ݒq�.U�l'ۤ�����	� $��9:��UL;n�8T撥?��^E/L��SO�Hݺuo`>� ��*�B��^�"L窎�WҁI�?�R%���p�66�^$r�x|ODg9?YQ(#%%�%�F�0#�Z��O�P@�]���J<N�U�,t����;�_��8��������
ЋV*�`ܾ������`�H���N qJ;MT@����7���"��}�`6���$&
U��%E*Y���[������-
�`7� Sj��  �³��+�g�f�&��;�wb�N�0����VL�1�^fMj2Q�Ɛ4pS�'&��5�"i47<�MMk�y<S���z���D�S��������"2������N6�U��	F�)qތ�9F�Ó� r�������~?�b���R����%�Y��Y�AS�9.<U���/2̐�<F��ӥ���Rj�Х�d|	�ǉ�%Y}��
Y��5�m8�~o�����m--/4;m�,�Ą��G���c�rFÐQT�B��y��!�;v�֨�P�{ۤFoY��tw,�ٮ�u�����zA�7iȶ�a���`'�4�1�ip)Z0��rh��p'z��~�%o[Z\�ENY�0�ؽK��Z��Fw+v�����(�p��Xù�4
-��B;�4�氒����Q@=�I\��ۏϝOრPeO1�b�@4����'y���}�{�^X������!eUt�
�9q���,+�.����|:s��3�<����?���O>�$O��6v:�,��od���W�8��Yb���y�)�=������������?ϻVy��~��j��0�QU���&WM���.2\��eW�9����@���[���;�ݝ�~��s��◿ĵ���������M;��9�K�A�QP�%�Dq�5�d��:�^(ɵ�:D�M���6�##�*kc��*e�O�W���RX}�?]�h�!?5���1Nh��י0NSx�"-ҡP&�<�(��>AP9���x}�����B��똰��U�Ĺ=�x���n,��q�Ɖ�e.E�Sѳ��a�Kh�,#�	ǩ��F��g�����$���D�?*J',ШQ!�x�an~^  �V4�f3裚��A�:�E��� �*�K���WH�NA����GE��]�@J���voS,J�+�Hs�1����42J��1I�V�w�Ν�}���A�7N��q�ybq�"M�0�J!Әo��F�x���(�3vR�}K�rzQ���x.�U���[k� g0��l�:n-c<w��h�ba�2B�{��Չe���
��N��� �]HVL�Y��)Y�[]���4 � [�K�-��p��MfU�BU۵� �pƂ_传<���0�j�����Kj/V;��s2��Q4و�% 9zT�-�r
� ���Ȗ-���B:!.��ƶ)�&�A[Ne&�;٪�G*�U���?�B��ʭ�-�L���V�5�!Y��y2��%�D�p��U��K����R�@��2���C����U�V�V��(�R�L�$��d.��ϝ�5�;����a[w�#j����Okf�\bB��-+�"��鞔�5��ؓ������������?�-o�R7�뇆�>����_���q���w�w��Vu� �fy�S�_߶-���$Uw6���\����'�Z��2=ǶB�ERJٚ��F�������=�F��������9~�	������%�аh�4Zh��
�,�Jǭ{n{��P���fu�tc��Tf`V�f���>Ɇ��_SP��E4�s�ST3�E�T�,��S��k�����c\��U0�!~�P�� ��	�"V/� ��(]cjɨ�mA��Td��T._T�]�VX����31K�4�7����>	���~J�d�wXFj�w1���Mdpy�@-@�H�ēD�3a�����U)�����ìP�W�df�V��RJҫ��"U�pF�ZC��ԑ�;77�������X��iu�a��Ȱ̠����7�oa�~�7�tgk��>������$F��لKg����"���v,ǧ���߿~��[��ba��]k6�a������-���vC�4V����������&1�{_X0KH�eL��I�&iRa�QEN��$�]\O&pUYӤ����C+B�;�/���ff�p��y?��OEal:�`d�M�RD'	���`�ĳ`x�#�?p�/��"P�W��Un�|h��9~�G�����?��?�����^{�iߪ�߼�9�ʭ���=[Q&��M$Y�%c	θ�f�Y.�^$T�����){I��p�V�~�_��ϯ?a�kQT[D�(9������^y�'��򗿌���c��Xø�D+
*"k֕f�GI��ݶ��x�˹��d �<fu��j�r��ÍK�l��Ы�S��?aE��S��?��
GS3��.�"�߷��1�Q�aY�?�l���](LS7��*���Y���Ri-��aQY�^9D}0�Yɧ�@Q;�%��9��ӏ�A6:͝u���;�2׃P/2�7�h��^i�v�sq;��B-��T�,m8��u�6F#`�����Z+O����z����DId����F�H����-(B�4%�R��T��FD':+bR\3�ƌ�@p'�j���>���k��$��4ҋ�C��0�#R�V�!�5ss�jT^��q �Uh�S3�6�N/�L������-g�k�%�֕~�Q/,���t0լH�4��ju֎0p?��:0ii�'�DWk�m!K�k����(�^��V�s��o~��蓮�)�I��(Y�ܦ����2�n�D�GH������µ�.~fk͎�m�N�S<�w߄6�XA-��{D̈_gwε2��=�\�0sb��X�m�K����f�V8��cʉ|fQ�F�A�s$Jn`�g�?夻�t�"I�l]-�H� {�����q�����̕>����wI��X�|	̪%{��$�A�)��ɴ?� }b��MB\�W���^5�,7E�q;�+�M�f�6���a�!O���/V�ȍ�'P��6-�^\Ұ���|�|���j3�e��8~^�L���v��$4�l�Qæ��qʴ�d��r�?@��y���n�;o����ϗ�5��oB^�A�U�e���Y��k_���eZ��5�s�R׺���m,��۾�Q�H�K�Ԉ������w:�7nn���U��L�lXz푇���#�u�a���~��78��8mʇ�������E�%L�(�����fZI�M$V��n�;�,��#��b9��h��=j�J�$��f�,:S8&�����YaU�|*�S*"6�k�qI|4NB۳���R���C��Q��7����h���M��j�h� ��U����}����
)�0p�`4�����69&f�A+E&o����-s�&Tp#YI>�H#6�Ua��<�=u@�H,�/EZ$Nd3�1~C���(�ݰ��������̨���i�$e�ǹB���6� �۪�t�+n4�_�E)!����VxfIX��Q��;}�����\-[s�������3_��>�O� H��Cc\�^�N�E,qf6�q����g�a�y�|����>:j���@���3��7�-�Ϝl�O���0ʔ?����7��7�jÈJ�͕<P�4�J�U���"e@�ЯG��u����}ֶ�s�U�ܫ�ݚY����ۻ7ڍ��꼀~��^�ѣi����{�����4����J��F�#?p݆��oj1���h����ܬ�B.���Ҥ�T�a+��S�{Y!�]�7�KJ�S��i�kX�)ּ/h�U�b#��Ft�
��-ϯi�25���۩W��8qv���4H�0>ah�c.--�w�}L����j5��ZYM��Q
I�(����M����\d3�'s|c���,�ǈ�:�*�����"Y$��2�'yo�_^�;��y��u�-uuuy4�ۖ�0�l�tt�P-ʆ;u�8��z�WL�F3�\M�s�?���R��ݐ�ÏXF���<�@�+��|�ȅ:���(ht��;x�y���bc��!��8���$� s��YY����$���	{Y���&V�F%b4c`(��.'R-|����F��ip��&@
"�RT�I��B�j���sgc�a������#���o���֝�O4�Q0d��(�.�V��Z
y��9op2;��:�q[vvv��3�����Û�677��ٳ��l<����p��o�� �<�U���GT�nS�
���a������eF�x����5��rT����Q#�e��+�Z���q8�������3���G�b�v�66�"3�6,��C4o�E�3*�_��m�c�����������DV�/�t>�|#SbJ�%!Ve�	��Ű?,Ŵ�"��0�����Q�3O�@]C7=7��Y�g����$63:D�,���8�7�˴Y�7�I��pF#���a"z.4Xo�����e'5�ejF��kN�Qs�{;�+�_�z��"s�l�T�RP��hNFpeee��k��(NXı�F�1��D-��,�TΩΓT)��ŨJ�Hf̊���PE�*g;r�vr�� �Vᛧ�*��1��<� 6�9�8��_�ዜ��q+{�K�RU�?�
��3��pI��(c�Z�I<-�Ne��T7��U=,�T-��띺��.ى��.gi�w�=�S%��d�K&f��,�g�OɁ+�pZ��:��e{Rֽz	�e�^��G�8��an��6��\���\A�.�T����D�i���vz��^o�����믿>���H��IO�(�z�ݽ�b�s��Ʌŕ8��UX%ͅo���[sN�>������X$�L�^E���7���;�n~���g>�8������P�4��9y�^�� �t{���_|KsZ|ɸ�tDQ<T�[�I {ue���K�p�b�tc�����B�KKO<�Xa1�D�`(�nm^�tynno���P�F�!�"���+�c�Â�ܮƲ��N��#D��l�=�����{p��4u����CD{��.ݔM�2$��(Nb�sk���1\H"��T=(�\#��C1����C�@�FԮHlz��)\ǆţ��A��$KT���$���I����&�w�$e�ȁ=Ve���H8Mm�L�`z-��wZ�t
������;{�q��*B��� N�q��8� K�b��,F��ͤ�iN|^a0�_ �	%��DY[��#mA��G�[{ݽ��變:.��G�G�?pf~���o{}}}iq��'j8���^o�O���̍CRB$2z��'׮]�j~��e1q�ь���s�V��K�������_���~�՜IcjA�XeӤ�N�V�i?.L���Sg>g[�������O}�3����0 z�1�tL��1� �cz�`�w�D,T��������z���{<�;���蓁�"������� ��%�O��dSST�I
D≌��/u|�MDv�"�X�y��/%j�J�tU�Dq��,d6;&�q��]L :l�8�S�ʓ)��1U��NN�n����e6�L n�$��b�ʍ����iB���YSn��m.�ފNtT��i������%B0�ȀI��RK���������.��~D���a*V!ÅT%��ғ$�W��#v��Zʠ�0�ʄ4�o�"౔�/��:��2�<=ʏ煉�;���$��(C���
w��4;{9>!�s�=�V֖�L^��%s��X�bg-��l�\��B�^������̠�Z�\��N��p�^�f��|��N�X��!7�^^Ђ��� 0C^()�jfc�`j	R����S��g�����I��Kv ~V�kˋ,Ѕ��uw��{E�ʥ��!ZL��f��6�o^酗<�z���k�]�K��^��,���2 �T{�u�����ēE�md��IOkM߫{�z��jZ���F3���9�(GP�
�_��ei^��Ĕ ƪ%_���
�5I}���EØT0v&��N�����:�A�����'�
��T��q<z�>̈́�6�v����D��4���V#!���E�J%5�('Qd⾤4m��������0�Qz���TM�$v_��6m �N��h$8��h���o�w�R��G!6���PE9`|9�$�Ғ8t��B�����nw��b4,�ܫ��z��}QrJIJJ��8jҚ���T�vNB5��6B�t؏E��^ !�.̿ZM���)8$'X�ʔ�C5�,;Y�����/!��(���E��yu���(OljOJ��1:��x�U�d��<�jc�1�NFݳn~X��`�`2�(;ű>�>l�V��R�"�V�`¸P}X�y�?�}��)��eڕ����Jm"y��|WW}��nV��d�SR�r��8�d����)2��X��G���o\�x���tu��)yD4A`��AZ?�������Q��f=Ž���4�#�q�GCJ	kD��
��w1��l.//��^�r���<���۽mj)b�Ǧ!lE>�7J������ޑ���iO��:@����S|套Y(.�֭[�F��ɓ@,W�^�/_��W�<|�뮻�4U�w�w��H^VQ66hgqqwq�a�4s8"�7֎����;�mw�Ԩ�f�a,x�}x5"��iܸq�s��]�O��ðtH�2�"����KU���e�j^���^�����KjĠR3��&������@�P��g( <�����lQ��P�'�oPU��0b�� �p��iKB#ʝѷd�
�x�:E8|�3[���޶�zp$U�'<M��
,E�H&���@�а�fb �"-/-\v�kk�3�G���~��{��u��fӘ�_�y������?y��++G���psk��xbkk��w���G�9<aGz�d��T�3�ݽ�z����CbxHR�4Yۚ�0;kQͮq��cgy����/D}�*4ܭ�f��1R�XS|�D�� a��@�A��&u͂3���#<;��ҜsFԭ���ƾc�gX� N�����|A�F<H)i/��5�D'�����&���I����$}D���}G����]B��eE%�"�j~�*E������5L�����V�PU��[����ն4Y�?, Zm4�"Wo��1�G �8�Ή*�D2%Zm��,�su�I��M	sa���!ܢ������j ��U�j����`������Q
�pJ}�(U�0J�����"U�*�FL(��W"1�,�8١ij��T���S-X8�Ͻ�[��l�9i×a�)�+줸	�Ga!٫i��p���{0e�N�h��D�gRݛ|����u�At�����¸Ɍ1���>�%2KD�WA�|"
��Ϝf�E����J��s��Ƶ�w� ���*��Ky�]��s��l��A�����`�Xɱ�K����P�����2!��XY�(nVJ��q��q����v;�յ�V�k���V@:�49M�	z�$9j���J����$^PkF0�%�Yo5j42��BXЊS�Wlo�7B~��:_��x����b<$�Ų,VX�a�sҙP������^1!�q�X��L3�3���ǚa��(�Q:ue�s��癁R� �o4�yo��/���4��p���~�;���������&V:*�[�5.�qRRE&+Ս���o���|ek��ݢ��P	B�,OK�ߥ�TS�,M�Y\�qZo�:��Ã���0��JAօ��!���	�Δ�k��+�w�WW�'U�*������<�~:E�$��ݜ��a�P������H�qlS�@�K͙)��jZ�:.%{����R7�B��'��72�Y�*���{�QU�R툐^��6�*��1N̳{�΃�}��MM�J��a|����rk7�s��N�_�<ʛ6Ea\e�V��"'��}���40i�&��'II��-wV()��ܶM҉�{�* H�U�3��L�6"��<�B�Ni�Q��<R�2��J�^�I/����{� K��J,�|��z�WWUo�F����J�H��U�QGG3�5E�m��_����a�(,�lO�g3�ES�"�$6 ݍЍ�j����r���}�vv�"�����f-������{���s��SSS�g���g �r,'4ǵ'��66���;��f'i������r�w�,�I!,rl��������Pt��^�s��u������,-^� ��W_R�dy��[�^w�"�q�D���w��uT�O�6��b�7g?��Yj�
话~�PM�D���#��؟���I��CP��{y�dS����RTM��#�R��R�Y��ĺ]�#��.��A����]���+����KS����m�-O��?��
g��P�ah���%*Ҡ����6�4HEv�$OȔ*�NF��M��9^���J�8L���~�ktq��z��JI�G��W|xFCbb��E'M�LDy�ʵ���l��/./�~05_\��*����\���_^^�����Zm���E�t���w�w�����0�ÄFiP�B~ey<�<H��5�l��Y��4v6� ����^`ydhsѮ�K%��~е3����i�_��x���q��Z]]��~������w��=Ǐ_\$����ʹ�o�p ������_y�����g>s�رь�p_5�����j c�fg�v[ͭ��(�x�i�s3�W�*{�� ����yw�rP4PLQq����m�.\�[�l�Io%d}�����M&o��*N�c�777qQ>�����C�m���a��#A��\����F|4N��>&	��%O��X__�5w%��˥Ѽ�t~ i�"����I��V�!��N/����G|0[�����ni�h�@}z� 1>\�.�uÞ��ؐn�mÔ��k�p2N������p"���;�e��~Ӏ�F�TS��ʲi���v���j��.9
��L���:�� ��I�X	��4ߕ��$4�wsG��>�*ț�,�~�onR-�{ t�����r!��mlCe`mC3%��u��ÚQ�!Q)����׷�_�W_{���='�=r�ݵ�h-�o��|>�)�ŌM�X^pX-�"��J�!��0�Q�����݂���i^ �$����$��B����O�y��>�Ⱦ}s�c�8�v��Ҥ�$�(�j��U�I�YF�m���PJnِy� �O
�B���G�Qr12�R\i�ߑQ$�>`�Ҕ1-��:C&��ըXD��~�� 	;��R��&f�j.ouJ4���#�|_e�P��*���� ��(��#g�O>O5��v��@]���$$<�/_	�uz]�L�m\����ŋ�)�:�
>HmJedh��i�ZU�F�zt�h�'"4�[�V�uFg3��M�I:99��'R�S$"�0s-;{����Jй�Ѻ����O�3��'|�����I7@i"�)_�3y=�nJW��� ���{�n�d8��������ǢL ����!�u<2o���f�%�'�f�����=H�.�矯����q�(����$+/�(P�AN�	u�	��tp�$c|����d�o'�S���8�9�pW<1����&pZ.?��.��W�O�R����㳚�&��驱0�Z��Yt��I�<�s��e[�Vke;�u���l!cX�_�YZl��7�m	��8ݍ�H�ZJ��A��p��6[Ol��4�z٦�O�㪩�G����� zC�]�x�\��M�b 
�c<F�Ѝz��1W늛�����ٝ��KV��Ҍ�]��ҥ@܃شZ�ગׯ��p�[:11v����OU��ۉ�"�KR��`Ue;J�$�Up�]X����M�L�J5�p��%�� ����+*����z���(�9�mt6��n{� �{��8��j^��l5���8㥵��\ �4#3M(�"�YnL�F�3�%��%Y� 6�<���r��1���8�k��7����ג��%�&J�ǫ�6$�����B-���ppY�`ލ��E�sմ	3��X���AR.V�D�5\�K��H�-
qU�a��5e�p5&`��nkye�ۃ�і�FGǽ������u�K�F����臯���ѣ��3���#���u6�uo~Ʊ��Y@��h����ޒ�)|�F� !��&$у��܂s�FUR08JC�d�SSڌ��
�W,V��Q��g��V��n$J��<'\���B��͍�_~�z�}�fnom��(ǝ�9s�����}	�.��X�9�<j9�F�X�?;O���{�5���<v���D(Y�(M�V~ܭe�5��(�Q���f���������"T�>����m�Ъr����e���\�ҡC���Z����(Wid�K��Ƞ�Q�β���<S��%�����_R��C�im�Z=Oo�j�(���ej�w�r����$�H�.�����,�$�$)�N�ZU�=5����\#�|��;9F:t�����.�������d�:_�p���I�'�z�>QXLc�b�̒��k,�9u�I��Q����T����b����L�u܊7�S˒ؤ�:R )�F��ka�e�iF����j�,�m6Z��xI���m(�U� ���
�JB5�#3�煽�R"_)�xc�0N�i�q�����;qbb�>2�)���ݚ��3fJ�����]H�E5�R�'���l�}K	�bW8�v�������~Wj�X����%���K�K�?<����t}�f�0���?�Z)G��S����B�,�%I�A
�����;�<�E�X�����́j�n8
�e�z�����q.�ph�f	'/�gLu��5�� RTK��4k��u���'���r0��6BեG����ЁJ�j�U]t�J���q\�읭]*�`#fu�J����[Y����
IR�$"`G���(��N	nD?��hR��&�,x���6�`�����z���iH��ȆXT��	�\q)�FϞ�x0t��Z�IS5�Vvv��g��@�r#��wx�m{~n󴈚'� �fVq^n�NZ
i1lO�$�g$ ݨ�)�~�}���		;O!��Q��@���g�3jQ��8��؃/Pc�RZ�\ 6fy`����x��P/�Af2Oxċ9����K����_��f>aQ��%� ���G�UR�,ǳYc������]������	�#=V��p��T�a!�� �n+��Z�@mdD��Lj���8�,2��6�|��}�F��
�ttb�9�C����H���7{a�l���U��5���v���8�h�)��ȍI�!-��� WLC����Vײ��7��#Nc�>�����.�}e�ɪ��a�<�eR$Erl���&������7l�d���me��gn3Ih[�����-����&����Q���0\�ݝf�s��Y.Vg���}ڄ[;=�� _I��զ�G@�p܆S��>���e��!<@>YN��	���2X�U��i?�į��mm��J����q�&�0࡭�U�t��J76�D4�N)�Q�Y�âl"n�2��d�Q2��sØ�i��HC=1,B�z?�t.�R�t)bJ�%t˖��g��<xpcc����w�������Ç���;JA>��jb.8��#�|e��qx6C�R-N֛�+�=�@�<�mu�5MO�����2�I�g�Wv��}��TE`�s�����*1�Ә�;=��e&[����T���/\���3�?G�I,���t�3���w��vu<�e�{_wL7��Q\�����.a�r ��g���C=433q���w�K\�A�,K��U��_�V:���U1/�v���JUa(jJ!,g�X��n�
���,6ؼ����/~�X[���ޖ�<��m)��ItA87�~ߨ>ʌ 2�#��D���N�gڪ9f�_ F{��=٫G�%�mt66wK���z���r����}_��:_*��}7q6�8���-,���<L:�	 w�OL�cl�<t~����"�2�X���[4�2�BFh��7 ��5�kNHb���t�����K� Q+q�ʠĚJ�+Y}
FS�5|��S�T��W�%���v��i��I���<kvR����`�Fی�\��+bا4���S*RTR"1���.��a��,W�z� ~�b,Q�mBz]��������!?� _���
������
���@hpU��Fja��Z{cm�nUJ#�)�E�qdeڞ�R�I�51T6�̇k7�]���%�U�c�֡?KsT��a(=i\�\�R}xsկ��v��GŔj�w�ӊ��5ʯ	�$���uۚ���&1u*�Z���h�������K��H��)��
��t�b��<K�Z�I��6�~ȏbSp� ��p3������X&�~���	�ܯ�H�ـ18�����B��;�~��h�<�`��|��@�|�M~�5�dDd��^�=9R��I�!�;��p�%�6�~2q����+y��d���ដP�����$�@*6�:˷T��@�g%rs2�2�pˏ�����)>���F>]NX�r/�G��)s|�x��O�����O�&mfLkf��	�|�._��#��W��*PƼJ҄	�<p�KCx��Fb:���_�Dc��ý˪a�ܹ��/_n��$�*yÂ��� R��j{�V�K���K�����,FP��������vgL7l�Ӽ�&*�a��Hʕ���ݽn���߹p������S���Mw`��R"}Mӯs�����CU���⹩�_AaTA��v��F��M
J���^SE�Nb��Ș*���c��B��{^�̉�9Ԧ�Ku� ^�N���r��s�\�����.�)���Dۥ"У��l�ʵ�C�p��6���HO�@�,~ǌR;������*�V*i����$v+
�J�iX�?��<�x0�+OUb��%�C>.V>!$�a���-��I�ص���蜂~*?.�x7L֛~��h@wث�E�_�=(��xs�h4cE)2X���0����3�*���j���ǭq��������sww�q�Z�<�  �Ʀ���b��5ЕH6�N���<r��� .)Օe�[��ڇ�����`�H)��b_����i�#�y��o���aS�dC���7���w�x��d���QE����D�t72R�vZ*�1T�1�,	��/��Tp�����f'��$KK���5k"2{J�w���г�H��*q6�[4W�[�:��)ʅ��=W�a^`I.^���$�^�B���W^y��_D4��O}���*�$���_��oΝ;�z�b�$����}��t S�8����	&!u�2$'��L���q�����yjw�,�τRf�%���O��y�a�ٙ�i� ��*����1���~pn|r�u��8�`��������m�,xE��aË2���^ղd*la�:M|
��4�üI�7"�S��G��8U���
�,F��iSEk�P�E�銘g��Az�x�����hF���i[c��QK��U���ͭ�@��-���Lbb��a�i��ic�C����è���#��������E,�W*�����M��>|pfzR�J8L�aԃ��ROU����:����Ƹ�8=���E�<E��eÕ�TU@�-F��W��|�����F}"�:1Q�� ��KF��#�z|�m��Nb����/�%��lIH%=�k��y:�l��)"�@а<%]���7��b�Je1��q�����$����&���}l�����ݯ��*&ŵ /�Xթ�6�{�:�pH�Zgu��T�d;7�CuoU�@��jm������U�WE�!�m�4ʘFΓ*�*���LF[$���ӠyK�E���,�ZW���P���S&=�Ӝew\7��U�P,�����z� ���N�[����BM��6���r��H*��q!��FE�+wR�����#Z=�y��b����x���(J\���2g�b�2�K�X~8� �|)��C!����S<�[��R��������r�`�������so��dr3O�ޝ�jd��9�l�H���؞�N��2b���(�6��\�ܦ|ww��	���k�Ȁc�������ƤZĈ$5;�2'R��3:�#�E��Ky��d?�#�op2|ɬ���[0�����؆j�KQ}��U� cE�B�P����QU0����v�ݵ��x�͡��vaA��-k�������6&r��BùS�TO
�w{���n��0�A�|��%S�'��~R��i 8@ǿ�G}��v��� �Q��a*F�1�
0� ei����D�u��nom���eE[[$�F��R��H�XP�%�:Z<�j1�s�"�%b�s�A�l|�(Zu�$�X`0_Z�g$����K�Z�W�MǊǺ���;���>��Z�X���$�X��,ʹ��-hcU�W>q�w���p-��o]��p�Pf��d�t�Z��-@{O�����x6��˩���:�/J*ud�Xϵ��k+;��a�+��Ov�v�ؖ*cf�zaq�[/�襷�l��	���uQ6��8Hv@wM#���c�ѭ�Tȓ��G������_��̶6�u�*�i��>��( C��ؽ,����{������b$���C�n����6��<�bi���g�l4Z���?�ɿ_������7�TB�V� Ŗ�C�p�I_I��p��Jw3���su�&�!��"�B���7�`���㙪U�'O����h~mmm|z��G��4�h/<˖Q�Qj�OG�W?�s?���/\�z	{�������X���n���Ø>�B?��������_p��F�{�A(�H���l�ǩT��쏳��z��Y�<�<to��2�@|̎�-?V�K_�ү�گь����=�NGx���|�M������y��P�$��vX��8\QY��J�2�̟�8�5��U��� 5v��~)v��eN��Z���Y#�7�V�2��:���s����`���w�Gp\�Wߧ����W����{�>s���l��$��hک),���e�ic1��?��<b���1�)�Ł:����`{�>����2� q%g��&r�~�(�#�u�G2U�u+Ʊc��c�Ħ峊���,}�]6���%��=w����(-�h�1��?����U���}���W^��7��{�GgSj������~Bm���hmzzrvv�����'?y��c�ܱ��~���ٟ=��K�K�Kْ4��O�����/~6�h�D�o�~'���!�ae����}gϾ�'�'��?���e�D.�w-%v��R��b��� �0��dq��^����H��Y)���X�W�w~�����c?P������9�kC�L�S-V���iNjC�z�v�����,��@ٵ�:�M�J��vm��mn_%�[�1����Q��x)���_���ciD��mѰq-I�n���p�u~�����j�F�'6"�XZ���aD���L�a~�ixJ�40�Ȉ ��{��2�X2�V�Va�V�����]�ܳ����^��il�ťj�2��O�"�k;��aO���̥a��1�<�,.��j�/�T��V�],��8)��0$�w{�yV�O�L7�-_YX�����x�pe��l:a��p���-�"��@����yp��k�,@�1�b��)�eljEN*9�Xs�f\('�1P>(�43?�2ZA�2���U|ɲ�RD�ă�~"*ҳ���$��3�Iq�*�N���vC��3���7a����`	]���1
��'Sr�8]J�,o�<�!+#Y�CR��Y|!R�)��s.�]8oi������3�����(J�#���D����������?�ЃضϿ�r�p6�zSU�h��J�>,�Jc�6>����7�<�t��e�t3�4�)9����O�v���+����,u�+8f�&��#ǵ}_�b����K�]]x�V��{�����7�O���|�����++��L���4K�SM��C	5���ZI�2�R��Å;�B�i�А�4��%1D3�-�"���XP��ȗ?��eC�ٽL�th������9�zKԄ�`�8��k.9�h�j�S��Fqpi��Ta{��}��~W%��Y�lY�������=�Q���L��WW���`������#_ɪ��`&
��!1{ЏG�D��s7���)]�6w���V,�-�Z�u} H��B������������~�ӯ�p~mgsdl�O�f�C�?&�6�u�1,�։��B��9���ݽ�Ε��ɑJ5����ۛ��׈
���Yl�f��,��*�H��?���8p`ttt^�Ly��B�F@:4��d{�h���heu#L�?��Ǐ��M���o|��}oeq�d9;���Rݶ����z٫��u#�v�#�I�F����_|�̫G���_�\�>	�����>�&��Cz�����t�6׮\>S�� ���y(30���X��U<)����С�V4i�^i���u��muY�}eiSه���0+�2��kQ(��7b�`����ƶO����@�b2]G��կ~��w�9q����9�N��� �
'�k<�/"�*�����C�666����u��渭����*^��=��OUD�q�o8B��Hm_ 0G�,������N���ܹ�i,!t��D��X��ݜ�ms'���pQ~Л����C�+������7�U�?��Ѝ�S��1jG��o����5���_z���@@2���}����q�Tj�� ���
���;Yp����y8Tt�ԩ/��w�}w�>"��p���$Q��κ�0��,AD�D{6`����z��E��W+�$b����߀`�����	4������G{�)T���OM�L���zFI4�*|䑏��/}���~��g������ �\���s���o�����Tju�R��h{�r�6���=���wc��ogϼ��@l��?�w~`m�0��)(��e^���~�!T�{샧N�|��򕯼��KZf6��`	I�'��I @�H;��Lol��3�i�?T:M��&�h�\���ž�s��q����߼ʬk?Y��B�ϸ���Q�T@�������|�2���܆E*�}2rT�o߾O~�3x�J��8J�S��  ���|�r?U�Sq��2���z:Ús�а�b)w|�-=Z,��H����q2�ڤ�d@���3��W�Tr]�o���q�>��f�͟š9���8bf����R:|����CxP���8*���
u�(e ,���[j.����4����waO#�-��|ڌ �
sj6?A�������jH�3��b�S�R�H� �H����w	��(�	�|��)Ġ�E�x�ׅ#0`���i�����ѽX7H˿dLŁC\i��J��&p�.�a����C1����k,zE%|��SGP���ie��ȯZ��ȱ���yl{c����?��p~�Ɇi<@[u�۳s��������g�Ւ�3�N��������w���r�Ŋw{A�HmDj�b>;r�0�_�؁���?�����G{��˗/7�[&�̘A�Ǫ�q�w ׾�N��"j��&�9^�)|��%0Xc�'m�o�ꖒ���j|w�^���jE�i�Q��ΰӄ+9G��S���v��i*�B}�225���"�<ҳ$p��^Ծi�� p�0����Jl����)��3���P�J�����Ѓ^�q��ٹ�n�3m=�	�i�[�"�^�����/�<��O,���g���O�~y��îf@�fz����a���gL��nln񃆽�yF����N�_��hxrZ�v�qH-�OL�2 �V��UvK��i������N?h6:��k%A7��$�-�1������ .���]o��Ճ�9����^}������?���k�����IھY��8��/,.,�4-,,<�bl�/ �4֏��%m�v��0��1T�k���>�������
���'��v/O��+a�f���`�}FP8ڏ~��ӧO����ZM}ͩ/<�<hK���Kf�����O�b�/��K��
�����'�Gs5?Q Ϭ�"!Y�/�a��{X�V������bj����W���"�������p9Qy�J�]X��^{��;���+�C	�̽L�\�qYq��]�|^|�E܂'�xG��_a�q�QT��a�)��> ��'O�D�;�h�G�ۮ�J�c�ε��J���5���7It꺁U�G����Dȴ[��|�k�SG�Uj�I�L�`�� 1�;�#�! ����ߘ���/���o=�0?U��>��_��'N��놺i ��--����@�Gُ����jr��'���O>���8}������~8�_ВbKQ��4���n���X�+����?�]�;���L#�~��b���U�n�����7�B��$�g�v�#e�����JF]��c�~{k`sK�r��g����!(+.� ���C=�M	'4�@�縜�l�X�zo�ݤFp��,��敥�!p�L�H�9�����$;_HT1����d�E�$i�2|$�B���;G�2cQN�a��"��JA�a��Ź�Q���,NI�r� �{#�{~%C Y�
8O|
p��� ����:��Ǡ\�b��5�/�au��h|��+�g+��I]���"3H +8g�^�1ӏ0�
|)����"�n��䛗DbN��{��$��i?��lp}�_�wJ��p|�^��M�>��h�������y��:x�7*C�iC�=m��Q��؄gfg�8N�Z�7�7������$�A �_w�����~�y�ރ��T��ݮ�X��c�4w���g��?���?R�����]2J��}>|�r���>V�cn�l�n����_��&71�k���(��������8�<�FU���b����ћ� ���-COjQ���z��յ����lwvJ�j�X��0�:������+���1�P�p���.P9�jӀT�ds���{�P2�h�n��4�Tͧ��Xz�f�fB�S�%�tAS�t3�+���Z��6�6U�-�v���S���BͫT>05���SW6�����������%��ӢF�ݾ�����F��W�}����<o��,��A�gz�����C�a5�V%J��iD:���ҋ�j1�z;3��z�D�j�V;j��-%�l�p&�n�kv� �N�ww�~����=x�c������=��;.>������k4vhN��N��ƾ?����u�_��_��x4�`>��S�=�����g~���'wvv
�b�+t���0oĝ.+:t���c�;����������:�zo���3{'�?�^�E�e�X���h�?~�����o���+�A��/�j��x�1����̾���,W�6AV9_�g>�h�����f�s�ҡ��<���ڞ�UYN�g���e��D��-��n��h<����g��q� �0��X>���vG�~�C  �_~�O��O���#`1��,��+��T�5`jL.�]�x�رc%���"?7ƖB�ʃe��qzC�F����ƛo�y��߹p�vi =�^	�	W��$rC҂$RXp����ӧ�[_]8��S������|��2Ƕ~�>��vc�}��g|����/�q�=A?v���v�s����?�&��aj�N��������z&_���_pF�7����
��sϾ���2����Qн���c~xbj�6�F�{��ۯ��:0'':q�gΜAD���z��M"��t7m�*By��c2ko�C���w/n��C�BP:��:绪8�ii�MEH��� �6��������y����W�I(hS}9VvO >���ߑ��9�'�2b���`��#^����Q��)Ѣ�>Q7�~Mm��O�'5��+��/N�u���q�+-p�g�����T����`�G�ZΖ�p�C�+q?�.ɸ��6-7� �8��.�\XR�ICbz��u���}.[q|ϡ?�x	� �A?m`9T��cJ��hyqH����p�I ���ppfB�ݕ�Wi����uA,�x���V�)����`ri�`������ Z����@���Dy����r����������s�2.l"~�3�������β� ,c��lll��=��@H�����d]o�t�����N�53�X�|��r�u���Z'�aZ��j鳟��(N��ċ]?>s��]Ǐ�F� ��ږa���qi��B��{���|�w6q>g�]���d�����{�BY��}�)nF���$��d�^[5Ҕ�������M]�z.h�8���A�h}�ӟ��?s`~��ե���S.�ퟟ��g�A��6S�Kc*�g�0���7�{NI��$k�P#�}S D`��a�#��%���
��,#�5�53V��O<�wS�(^��n�\��[Y�Y��`жkZ�c�\����M*�������_p��Vi� N�X?w�n���[lllbr
�s�ٝ?8�{𿯮o\�C�Ix*=��� O|��r�{����q��'/H��qq�Q�7v;��}�����=�(�Q��;{��W�}i{sk��v)�`��X�SߩW�+K=�S�ܙ�������<��3�Ͼ�ƙ^x��������.N	�\�V�^]�r���N�7>A�;�٩{O��Mw��2ۡN`�^F1:U�����}�#?�s�n�^������}�+_��իW��Ϫ�U^�sx8�tS$3Фݎ[�٠�� k�R�_��^{muu��9>>��祺��l�UG{���6��K�8?�7�y ��#�(����b<,j�7j��#�Ìݳ����;��[fαJ���R_X��d�j�G�{[I�qW!�����2�ܻ;33���⯜�cb�͠oY%U�� T�W5��\Ϸ��m���>x� n�W(�O$�@�{���9�)��C��35��XvFZUa�:���cv{�g�y��矉��6�&���aU�y���V���8k�:��o���������0ӵr�7~����z�!&na����c�~�՗�.����V���iX;;�7޺����?~�k_kw�~�7=5�?��_���?��<�{�9y���7�x#Ӱh�g�}����T�;�'�����?��/���WΜ}��'������kk��ߘ$Bt\�PW�K�(a����䖇��|���t�߆�n+!�ŷ�T�� &�5gr��]���.<�l� ]�9fQ���<Rq��K����,<��ŒE�y�]Z[n���A툋ڬC�gX%����l�fPQ��ǣp�8~F�p���c'���0<��a+��0m�S��iƩ/�}B�bw���3�O&OR��"|�K"�0�0���R8_�鲟E.���.����q	X���e^���	��8���/���yep���i���$�D�k"N�&L+.�[\>�G�p�=%v�0��pR�]���=3��K藼 �?dR�t1	kB
bҧ$k���ޗ�7�n����4�*⬧3T9ӆ�($j�ϕ���d���J���۱�X�Ix�����U�f����=�pgبtz�*W6��kv���~���"�M�_��g�8]��w:p�Ё�j6�|�?���M��]<�*x&-g��R؛�ǽ"U_��β���Zݾ�[	��6Ʒq{fD����Y�?Q�sHhE3T:��i씪#���_�~�g���=��=r�	�z[Y'�7�텘4�5�+"j	��0/���'�K��qC������\�����z� �j�]���~m�!JR�I�1�S%k�FO����kD<ҍ����Z�j^jf�~g�Rͬt�߭���?0��i��rJ#��lf�4����nR�}+�+����Y�K+@=���553���eZ�%�e_ *�RD*��7j��@̛�4J+PM�THKh�D��h���0�:t���N�hY����U����׿��ę�Z�B�!�h��jI45=��#(�����r���}��{�ԅΜ9��w�ܬk[̃�M����ꫯmnn,-���ؤ�l�>�0"]V"��I�a�9�|�����c�ҕ�����>s������
�򟺡���L�ofȯ�hf0�`�1׈`��𧭭-�6����߉�	��w�;0T��I�Tl0�� �Z$���6O���e^5N�*e���oMWaU����蚈8��m�b��V7/(*�)	�c_̍[���ܷo�5n��Kވ�A$��ҰV0����LZ�E�ra����8R
��u�~ $0���'���3�s9SC�T2���R�Q89!�4�^ !��m۽v�F0B���,˲繻V�͉k��ga�F���>� nuz�Ͽs��b����ُ�����w����#'�w{�Ridv~�����n�Ԭb�Kb���K/���sϽ����˴���~�w~�ܹ���[����ۅ���M����D"�v�ѳkH��4i�vqk�..--��ސ,��ᐜU�ޫ���}D�s���푨��P�����+F�(U9u��n��w	���Jio #�V�`��<���bA7u\`��Nf7�z�>���099�k��X�t��%��,�=�� x4���E����A��L'&�MWk���<``�Հ��!e������M[�p��(g�Y�J�+��M�oc���gggEW�Q~�jR��Ƽ&F\\
�>!���>+�L0���X]]E�we@��p?�β탃g�����Xsɹ
{�M!��)��(� |�cr�����:~�������`�077����(�0���_ò9|���I�o7/ɰ<^��̌gg�ē��=	,�ν@\&b?�O�)��*����� {;i��s+S�e������	ɮ��a|L��}v����W�� ��J�^�˧Z�*\��Ƨ�M*�R���������0
�hjr�;�pcmsrl�I��H�>��X���9qg�IGj�ږ��vyem��L�6�n��}#�
U��n���1�B��F�,�-���b�+D~tS� �+�h��`��?:�����+��z�iZ.{jR5�b��jo��x����c'��8j��T���������*��b�N=����b��ԡ�?�jZ��S=��t`�u�A ;<�52��B��9�M��?׊��n&+���)�	�r�jbc$�����̒���vͰ�]�t=ʀ�*��B:d��='7}��O|��]��tӑj��ݙ������Ϛ�9�r��Y�,�+�N� ��݌8w e- I�H#��v��L'S�ܚ~?�zxKNij�W��#:��0 ������҂S.���I�X�.\]����y�#G�X0ٸ��393���}����f�KȥZ<�x��EA�[h�v5D���j79���I�F�+U��f8�=���Q�0�5��ڣvc�y���qVlr�"q�.n��>L6YLQ�ųau�i�G�m��V����͞�h��{�4E	CБH�
�H�l�B�W��$�G���;8���C-���D�}";$�U��|\;�;��)�p��Y�\k����L4����������'zv��G��
�cCbI����n�,���"��h�HE�H�\�HJ�q��A�#m��M�e�CI����!*i�vΜ9s��e�FZ��3>V����~���3�^2L�Q�.�4Z��cM�Օ�����）�i�[!��+������[o�����V����(Ë,��Ơ�� i��~������Q�\�6�ڴ�Tm�TJ�7p�~"��<����#��9i
��9����{���he�X)���K��+
��.)s��J��X�I�t�Y(�90=B��5��!;���	�d\������aSpd8f|q"�y�ds�+�T�th��k˱aJ�j��2i��+�;�q#��S�i��-����0lv�)\�aC�,� ���78%��YI�)��p2�L8&���GNȉR#��H>��i�q�[k�'�d�:�i񅰳 �y�Z)\�k�s�yYL*�99��◱�_ ��8�ɨ���\�b��C���7���D�\�/�h �o|gyK��2��O�o.g��������H8,ch$�C�d$7���f�	#j��ك�]��|�l�O���K�r�ZL�T�G��:x��=��C�"�+�JʛMS�L^��VD��'�;]˫O��َܬXF`]���~/Lһl��cG���h�I�4� Jl�$�����{.)m��A������7��"���^�t��U�Z�p��O�~���%*H�߇!�.�p�}AA<�UW��2�ͧ��겑�w��ĩ��Z����8����K����f�zmD7�ݣ�����p,W����Š�!3����D��q��j)J���j��j+��ۡ`D7s�u�L��^�;6�L�J�^����Iܒk�>�N�`���
�=����1m3�\g\U`�r����X^[\Y\i6[��L�͌�F�W�[�Ne�c��trIj)F���2��JC�/?�M�	W'��a�tX`N �4�v���W�ҋ3����,mae{��)�<�����t��(n�8Th�X0���	�`c3�U���7��`~a���p��FS�=vv��V��u�0_4���}�EH�7�4s<�p���"v��1٤��	M�&euM��?�'���i�W8�yX"f���e�)4�s���^㣱��7�H�&�v˙� �n����[� ���q9����y�ȼ8�L�����a�622��x!ͥ2�Zx{:<�NAp�LS&����Q�a�QN ��,;v(�"d-D;�7�IB��Ë*?��{��+�4�f�`RO3��\���N\4�n��HՈ��h��F�1U��?)�:z�n��
�)�J@�Tv�/�$t\�e0$�o	̏NT�V��
vak}#��J#�~?r��fk�+k���y��C��Ԋz���������!V>x�~��u͍�����b��$IT�r0�eN���&FM+����B�Iw�-uCY'6F��{,p�~��N�z�~<b_��P��#p���<�[�d跨Dݢ�H�w�Ci��N���;�vX"uc��"H}E��z��^����b�7333==������&A� ���/pnn/���`�IwA�Y�+�2~P�@񮹚�f��E�L�1�JF�����+W��<8�` '�Gݱ���������a=s��,�V�ss<�ylai���:��1��P���ɳ�br[U����_�s��Qc��%������GH�?�`��k�p¬��;�8<І�Bsn��Z����?�<n��b������v��¿\������8A:hE>[4��r��,R�������9Ra8ͷ^��D1��(��X�6�vܓ&�W�!d��e(FJ2��W����U�5�f>=^���w,��8Mx$"��;u>jc[㙈C�=83-���%�3�����[�������v�D@AZ7[;�qn��#���
�7�zkkg;�>X�mc�m�E������v��w�MmgX��ivK^g~n��|銞�R���i7����N>�͑��Pk���ږ��ql7D&^��짅�p��H˒d�ظ5��w�597W��в�s���O�^�z���pa��E͊��gZg�	R�-zO]>��LA���Ti�Cg4Y��)()�.2�z�Wi����5��b�f���,*�YH���>f�-"��鴌��*�)���mw�%����I�MzA��>��_z�{�^���k�쯏�K��:.�km`��>�36 ��S5�p�O n^
��/�U�z�hH���c�L+� �������V�9�C܋v7���Օ�b��ՌAC�1�&Q���T��l��.K�+%q�j&���!������z�D��|�M�.��B���c{���~������\�����6�^�����M M)`k�}�ʥ7�|���oY�!qK����v˭�o*}&U�Z�L�'�婧��ʹj��b8�Pʨ:FA,�*���;��9i%�by��/H$�DꀝZ�H(�ha�%8'Ѕm����2xd���>Oɲ�#.��R�@N)7*P��|z>=��GC�o�E�[�.���"��bƄ6�~5�pi��W(��2t�d�s�2���0���T?U�pi9'�1!AQ�3&8�����I�(=��v�@����Ɠ��@�I3Y�K�T���v���T����a��|xi�-v�����|�ɃwGHG�<�[�� �Z^^��\�:���;���#�м��)G�=�������R�&a���$w�mnm��f��R��k�g����"��IQ�C�{�D���u�K{��ٷ�u���İ��(T�:��X��7;yp�t�mfZZ���'��_seiU��:�^�d�:���F�`�,-�V�,���Ȣ���ý�u�	9q��z��c��}�r���Z��6��	D��f���2?K���n;�u�E��P��q�ݴ\ggk�ھ�i�-�w�v;[���G�u=�a�:����N�5NJ�#Dg�m�?�B4Q���^��m4=Ӯ���!ҝ��ǅ�~R����U����A�G�.)�5���� ��Ҙ�Z��ۺ��29>����(�~wD��F���M�*�*�nf�Q���W���F*��;�9�f+�mk��u�L*���S���TJJ�ޫ�h����&K�F���,>������^����79Z����� �
�6�n'��@�բ��F���TJ#���	:�F�Qb8�|^b(��ʍS�D�L����|H,N�qmQ��A���k��/3�!.�'LD������ES�Q>�=_�	d���]�3��5�ۺ��k��T�P�}_'?��f��28ס\"�Z�h莊;q>�@�U�, 8�*x��H	@��T3���l���J�6�`0g��(I�Bǭ��v�j�fw�z��i�P�@����Jb��ȔiU���i)���p/ :Bq4���X��_~��r�`��[��v�;��������G;���#/\y�4�6���Q�7�MSV�|�U���EiD\�n������b�R�0A�ơe��?��A~�P�fQ'h�_�5�$6,����&�D�F^X�Ŗ�Ц0�q4�Ӧ��@��F��C`��6��UF�F�\~�#��y`��b�����Ak2)��A��n��ǝ��899���-z�9}����'�dq������.^���G���As1�S���j�Zd`�����iq��t�4��\����N�cdNAwMk���l�傧'z���Zf��g���ȢA�sM ��v�T��������f�fJ)���c$��Ѩ��O
�.>L7�{�TOR���uj����e-x{�R�ʕH��Ǜ����O����,��x��@،˪�p6%I_j�2�))<	I%�U��T*;�"l�c���7����٤�P��	��}��~�������+���W�O�4/ӫ�W�y��'�p�\�hi�Fq[j�L��땨�*ĭ�}�"�`�E���NPb��P�v�b��51Y�M����l��~��L�j���z��b�~�c�o�l[�ţ��^U6�q��ե�il�8�����o����v�^n60J���Ԕ�O\V������9#�C���l$�G��l�~��S���~�W� P��8�;gj�S�+���Űݣ�8�XZ��m��Qr'	��`g]�!�m�o�T%+�j=�D�ENl��"?��v����#�KE���p���e2��W2W�!� �NAX'��)W��������9QOJb)$_){�0�C��t��c6�tF�Ql�8�~M���ݠeZNFnAr���:�����\ֆ����@t)�i�Ք�̠���Ee*�x���w)ެ*p]��Si7M�^W�Z�/6��Vx��w�����(1�.5�U���mOZƈG�FGf.]��{��ǖ��ݿ��Ց�^��o��Ct{{��S��� �p��׿�o��n/ ey#̒�XrT�B�[�:.�l�26YuM��L��juD]l��x�8%��j`��)��5�?��P~3{_��O�GH������o�X(�2k6�ܿ�����^�V�9r�����>��^���.��js�:]�4t?�6��csc�2Eap��%�
.�A�4�FA3>���NNNry�)���ۍ]�G�f���f0����ݝ���f:1s����z����N�u$(����������@�7�}��ޡVH�����o�F�F��e��.�i6�v����ώW*$a��xW�;8`I��GH�:a��۫<�&xk�������YX[����A�&?�Akc ��d�Z�Z����D=-�����զ��������ZJ�P07���AD�W�~���C-,^��'Í7)��6�8� ��8겇@���xP�zL��5PH7���r�RqK����2)�
��ib&)�0� ͒��5�-�6�d`�x}�w��$�\'���|�VL�U�qSB%��Ю�k�_��_i1����qJ�j)��D���v����~7�����2]S,za��Pe��NM��u�ʕ�om�4���߶���K�ݍjy��{��b�vo�!��5\z���1+!0�/�*�1�͈�*�-,,���C�?����z�y��`�c��pxY��וV�@׀�}����h�Y]t�i�4���)�
�@lO]AJ�X�4_:�#I�G-=�P�]t迂��I!#6�j�=	?M+ƉP۴dfR�ՠ�oH#&)XIU�tm�#��F�ߞ#'DD�� �?��ш����\d����#GLw�f	�4��]-\�n����П�~J�
�l�2]-�}���W	�s�}�",�up����6���Ḇ��b�Q��)��xF�o$��3)��aI~&�aC��$e֍j�(�sѣZ�Zj�6"ēw�h�n/\��j˝v��h���P��FN����͏�y�w��c�>��'rHC�k&��ai�!&�(z�_ s�TSU�g�S�u5@Ƥ��,@G������|m��\i����*��ѣG�bu�CS3� �@��v+U��DSB�r�� �ffgu��1�1u�� G'�s<qX��vRNa��5��:T��t��'5���n��Ēi��`��Q�C� ,��[`��J�h�c����S�$��M���*��:����L�`m	��̏�T���d���3���a� !�	�[�!�����oh7(��'���� �
aO1TQ:
h��rzx'&�'P(���t
B���1��2<��d��	���� ,Pi�����P[�%��̡b�'c�n����(?)�MB6�8��2�{G�0O�N��:r�Cx�R��v[=?�J%���ե�������җ���'s�������m�v�������_~�677B�^�����~�/ۆ���{ ҫt���""c�~F�?Ձ����7_���38[�o�g�g��`)h��a����g�}��g���QD\�0�٥��)xxw��V��S<ojjB��
�c��e6U�J�6R/��(���'X�7�&)�+U �X�c���i�vF���m��d�����c3��H-�Ɇ߈����*�e�9�S��N���m���kR����^V���$`�F|���	R����ja%�iJ^�K�q���ӆ�x8T�-1�Az1񧹹9hֹ��*k�d��E�̄s�2ܛ[ۜ3T(�Vġb��]7��)m8��� %���0��
�jGŌ��qx/f����L���}�˗/^�po�뮻<�{t����+�t���pl����m V�����O\^^~�Gg\�����;�q�+�O�^Y^+��M�̋�]@�Wd�.2q�L*�� ���F8�����	�=::ʂ�8S�j�/s�q���&aЏq���s�T/�/�� E~Agj�F��ng�z�+��Q2�q�=c2����et#��j����F���z��E��:�m6��<%x��~������ހ�ӡ�Wa�.�X?K�Kelt�Z�'a�\��7�զ8�'�7����-9���aSH��z<�竘KF��q/J�вibNG&N�1݌2|c)��(J��f+��~�򽡞�B)�C�'�d�Ylz�	�O��:LS�Ji�:.��|��l�����U�姲\��_91�WW�f�
܅ūW�\�J^��L�*pbQb�Xq��7�L����Zz��28�[�,�h�m�S� �������Ue KB�(*-\+�t�t�J��5n�"G&��D�F#��%��R�u�\�iu�O#��^H�.Uc�LʨbI��g�l�a��jk�v�Iil j�yl�x�w�Okml	����R���:����f{ ���8=���ۨ�]�T���CҨ�U"4��:��H�)6�`E*R�9N"r1G֔�6�u������c����'Μ9����/Sj.�����0�0w���q[��9T�|�����B�AhΣc"������9t���Ų=0,�[�z )@ֿ�o(x�M��)�ΑC�����j����F��Z�LP`�ȥ	\uA�����amm��"5�H=8R�I��NH1���8ʗ �jl��L��5H���7��R��c�\����i>̋��M����h��ݑ�䧖{�BLm/�� �y�r%��@p��#�����ոb%���O�!�GT�&��U�w	 �r���m�-�T{�ύل�����P�xPUdx��R��:�o����U���ssx"�ʯ������p�b���[�Ͽu�|�i��3��_���8�}�g�>q"R��(6/��m�G�����������˷�>��*�68O����5����:IJ�4ͯ����_@k�=�����K;<�j8 C	� �L��h�Cl։�������;�!y_?��m²9r�2��W����fpjy{wgؗO�T�r8�����_�������y��?��pČw��N��O������5��t���g��*Sxgg��=�O�S�q|�*.92�!���s�[[N�T�j�
lmw��T	Ƭ�mP�����UKncttR���0�mggK&,���G���2] s'�_s��� �>�CU�HR��>;� ��@2�/�&�4��&QǴ��x1|�*U��r�܏�
V3ǚ��v���M�Ь�qGBwPc�t�S*8$�gYI����1.�K	�l dS�i�T.c��1×��G9��9�LL�h�yq�k�q��9k�* T�fn�b�<k$0����0%Nsr֖ձ("�|��)�y����%Sm��������*山:�g,Ǫw������Vk$������w�u\7к�Sx�G����;�|3�2����9�Vr8�̮�∣�FҨjQ��|���H�U(2�b��D]drk�%Ա�9�[:&bii ~:�~���Qÿ�̌D�4�S1,FƝB4a�i�)�l��	6�S(8�"� �8����(�^��K]�P��Q�� V!�Ψ�[�u�l�����r%��Ht$���C��n�}uueffJ��p�:!�2�T�>\u&芴�� <��)5��x�ߙ���E��n��Z�J)�`?(�E�,���"P�Râ�A��Th��:�]������.��Dy� KJ4u�B�M�X,#�����I� ���lp�8C۰������B}j�>�k��p~~�[o����%����Un���M�y=Y�e����X"��!�Ȩ22��=�� J�wvcΎY����QL��CD�`�KId�[�aЎ�'�&���B��&� ���t9:q��EO�~��'�A��sM�:M����q�q~@�LK�o٠�F�G�8�e�@�Za�ҕ	;ص�*�|ـ@�\	��|J���M�/���<�=E^�Haw?x��7�x�Q�>���R	���'x�������ɿ$q�Z��d����$�l>6�n�V���'���֧g�aA��i�Yi`yn�a�a��Jt.��=���p:T�d%�����V�}KG��)�{�:�ʜ	�@.PN�-Lr>0��{o%�Y�	�}�=3"�����hI`�����n���}�ǧ�����?������������m��1��B,�$(UI%�jͬ\#��������ވ[�,	lL��EVVč{����}�wy��x�$Τ��Q=��H�0��O$*r�#�n�e���9n_��S��dD�8�r���Fű�����qs}�:4���' �-�R��f|RU�����s�յ�Kb(R;z��S�Μ9��f�՟��t���˃�"�"F�h.\�������o�����rbbzz����ŹBQ���_��_��?������n�V,���#`�j5��o����pD7D�?2�a�����f�7�����p�	�=r�[��g��������{%��?���}��Bmf�0�H��F\����'��-j
�w�W!WHP�ܸO?��N}.�(�g�AL��Zh�d]�8e�E
Ge�A��M�!��w
��Ϣ���%!�(	��+\�v�Qg�=�����}Hjzq[V~r�i��Jq�d��q����ҁ�M�.�Mv��ɯ�;.E%y״턳t�>]��/����W�47������0�A�I4c*�#�S����2��p���԰1�r��ґ�PK���lg"3�zN-�*lAr�,�'��s�$M�K2+�9�':ܔ��6��}��^dx���}���������7b��e��I�c�❁h1sxn��8فfٷ���(���e�|�۽����EI�p=��,�e�1�웾p��$��#�K5���/ؕ^���/P�CL\A�׮��C*��B�@�ʈ���xRx��\��-�I��ry1)����˚�J�̬P8Nϯ"�	��D!U�-�� �{��#�er$A�&��gj9�M�-���UU"���(�8�aP�=��vV�#V�����\���l`ܦ�c���+�>vpB�'SM�4�J�dm��H&E5Y7�r.�$=����+Ej�OCl���T/UpS`�,חZF��ᰀ���Vq�5��V���e�4#o�*�S��5�z.Q<A���K� �u��N嘇�(LqV)12I���Dʀ���~��7Q�	�D�/���^9V�l��[U�P`�ƣ���4 �K�I"l�V�I�Hե��B#E�[�ئJU� ��x�PL�S�a
#h3�Eƙ�'�
���:|��!������;�;�A'Z¼8<�ĸ*��@�)+Ul氨
�;�[�88�����T$�9o�#��5����D�Ϟ�j
8,�f[&��D?u���[�q^1*�o֟=��K/������'����V}kcc_�e�B�P���_#2�BNh�n�Y��2�t�2��q��܌�Z~�DX&��)?���s���5�qCVY����"���Z"��E>UN9�c�̤g�+I��b��[x���.#�7@X���b�9o�)s`�&��;KK�:|��!�B����{�9NVf�}���8�?_W&�pksoF1���]��i�(lQ�L*	}R"����iYǎ-9�I��  �-�a*��8����~��^�t0h�^����ݝ���+����R����|��w���O�>'L��G?�a��������ߡ$������p���tڑ���X�-j�IbѿȌ���S,#����9n�z��:wC���.)�vvv�x�	ز����~���Q��wܡ����rL���OEd��VB��2;-E��'d)h`��B�IT0�RL�jFԳ�Ұ�[!JcM��!�G��(�膑PY���G�u��� �?Ն�愫��gJ���T��,BFM�T:N[�hD�2� �Z��%ȩ�Mr��4��8$���J� 3�Xi膦SR<��6$�FV�Y�̞\�p'���5Jg�B<�� ��_#v����CAH�w|���8<WZ2�U�:��@���e?M�����g�
�܋6��TЀ�̴<L�!�-r�G�R�	 ͌m��	�E]�j�L����|��h�.E��(K��|ΊV��tQ��#�m�D`<�S��B�E����`3E6#ryZ"����2+�H����
�|1sB�M)� [�(��ǉJ3�D���2�q�h�F�ds O+V�d�5l����Ӊ�"L��px��|a���^i�uS��q�������*��n��4pG�<d��GR�����7Vez�d����lz"��iK2mz�)9O�e�|x'n�!&x�U�_�9z`e���ו�PƆ�{��A�-'!�#I�Ä�P"&p跖]|���[Y�%f��	!	�$]����dQ
9
�q�&����B�Y�Y@w��*�@:v��ԝ^Eհj�"�TP7ubo)]��ٔ��Z���e�Z#z#]K[���e<ISG�؅��[�4v�`��S�\�����ͦM,-��qJ�,�� >������eS���DŒ:+�+�r�W��Ɖ����>��X%�Q)ON��,�J����5�s�T����
��~gmmmks]��3	��x��uT�}O�t�o� �GA��H�cIY�X�R q���:��O�kⰀ.�������q
��>vLGJJ�ZBy��^�=l��5����,�@��K��8B|�mÈ�,�e�g큛������r|�fr��)\�PdNf�����)��8g`|�aWK�C�M3�Vd�D�
TÍqg�����Çz�!\0ϩS���m����c�e^�z��l���I7�(��8�_ "�n����C!b���P��dImuڗ.]b~��i*+a)��4+��f}�0�Uɦ}`p�66ku�8$��d�%F<��Y��ͼe�%~�8��-� �t;�n�	?�P�E���9	�$i}c��j�+����ٌ˔�$�I533�s���w�s��驩���bx���?��?��g?���a9P���օ�e����U �Ѳ���}w� _�Er�����w���)A��Ӡ*  %GX%Y��=�ő4�����_��_�޸�h�|��m��v��|gcckm�����3���ݿ���Ė�8.V�]�z�����(i���c��A̍sR���R8s���E���A���ʨ9�3�SF">���l����G?|�=�LMU)�#d�l�?�DEQ@�&�����c�2��YyFӇ�k�d����C?�i�=�qUtp�z=2��6���J�qA�O��h3�6~6,KD�	5�IJL�'�>n�o�i !�h��G�ؒOf�^J�P�pF
�FƮ�v�i����*/KNs�,�J�����@�89n�"�f��!�뇙>7s*f��t�DUZ{����?b�A�����p�V"��M����%����4l��]�+b7�6*�ڰ;<���I�A&D���З��9�A���=lw�G�[� &�7��(���2��Ex^�YdD�7�TR��	���ͺ3�D��BEW�R����ɫ��Y�Ax>U�
�2�u[�-?���P�V�oI�ʰ�E��x�	����Sil��mV*��;�>Voj���A:tI,K
p}{�����]���c��@8�6r$�4�J��Q K���eY������p'�1BQ��!�Q$i@�؍�|!�,�BI����EK�v572�!�����j�TO�|_Oa@dc�B�D	N\�N�l�*;N�ƹ�v����L�q,�� �$�Iq��X�&\�vӠ�7���#�K3\_𒩒ۧ�K�ES�`3E�(��k!�i�`�_Q��g��Q���UtV��=�e:9^SnRL�0ׯ_���>��3��Q�t:뫍�8G����Yy�����ڔ�xn}k�뗮��D}V�Ϝ>�LL覕:�ƍ�Xҩ�Cs���U���fk���K�V7���N���;uVL���T�]P��P%p8 ��sG�"�d�)�lvVWW�g��s�*�l�;�L�dc���/t�-�n<0�^�s�4$j�xi1�� a��l��@��-%&lQ��ܠDC���Ԟ�I�_e��a��k��~����@�ߋ��8��ib��8ǹ��_bC2�q\��e���s+�t
���!I�p%ND֌��;�a���A6�����4�����:K�1d��,�ͦ��`��hE����,��kd>���\����3��w߻��nz��j�X��Mo������s����ӵ����j�
w��SO}�_�?����{I=N�S�8�b������W��l~<�T,&���Y��և�@9"�K�ڍ׈��91ǀ��:{e΅+��^yF�ui����Pu�9S#������̃�'Y�����xwgs+��U��
���y�ر�~�]�>Z�[�|X��X=��g�y��Z���O�c3�ފիX#�{�X����h�+k���,��Ð�����MT�~��v������fg����łm�0��+��>��>���_�G+���:�0�AD�9������)� ����/���{>��U�U;g7]|���0���f���{z���y N\��P_\"���:zcF����L[�s~�$Xq��j�(���]�t���d�(l��,����{|t�:��-,��!<xq:$��Ycz�i�3뺰d�e
N���Ж�o�6�y��tzQ�ZD��N7��d����<,�e���|S�d��|���	&�dI
م��*+�9MWy�1���l��#gg ��8�=
��Q�+p���Q*RP��e��w�!�hp�0�X�N�J��1�+�������pnx3k"ᘤ�*8�q>������(���n�r�C56��=¥Q�^Suvo=!�ʁ�4亡;s�K���eJ�bͩ�������!��v;.�F�j5��tiq��	0�e�x���su�f��<������Y�z���Y�XȲ��(�>x��K�$�$f�Ds� �,��+������)�?�
{@O�BES-b�2n%��:�k>���I��;Q�����������y�6\�	�D��g�}��z���FF|�|*�"b�
B�,6jM�o�عa@ W����p&���F$�L�������AC3��6�<��a����]�5o4���#GH޷I?�j�8淾�������r�Z�X����������Q۶v����>�f��,�;sS"L�_+��r��&֓H����M|#�w��mv;����R�\��R��7�~������E�������f E���!Lq�#�.��dٴ�h�dQbf�$��"OI���i��� ��5���Jj��He�.-/G��`�n�TU|Q�����t���Gr�F�y�'�bZ����iɌ#���^)��z.�Ф��Ns�em�wr�܏�5<*W.,�ѧ�R��D�&&�������!g6b�'���x Ug�5�Ł�k��(�B@�{��qF/^@N^���l�m|F�OSP�$�������x�ej*7��P_[v1	L�Lc�>P��0�$pRcK�ʊ�r�Z ��|��#VXʌm&m��n<�NvF�� ��T����EA��!3'
�1����X]�z����&'D��]�i������v�G�<��#���4����3G}��#� x`�L�q���j��u ��'O�T%�2zTB7ͻ�箻�ƿ��SR<����qx6�pN�>���]X��?�4	H$_#K=��؍7~����_�2�_�l��́�����夲�L��I�g> ���Y�(kb��s���"mƠ�}v��9.�����0��?��{��:�4@�/���n���������Ϳ��O��O��/�"|bW� �'WҀ0{�1��x�}�1���˗/g²��B֌��G�]�J#g�XX	O	c�����[�Y_-��J�k���Z�M?~��#��_�����߮�^���;}�я}����a�ǚ����](�R굻�r��o���b��|���sϿ����D�(������x����N�9�8��W$-�4Ш���
b�8>rJ���M�n�b��?dy��7���f���1?$�拧N�X�Ç����<��WW������V�ؤ\ 
���VGt���՚f���m����d��MKѩ�@l��u��#j:'�)�)&T��Q�B��p�㰶Ic��tʑ���~L���c.�W4E���t��j+www{gGV��e���ĩGJ'�p�L_F�:1��E9S��8D���w��_���R�ƕ P� �V(�TQ�ߡ���4���2�$�MѕΎ3�~��L����w�tZ�n�F�=�����v���f��pn���!S0$(䂎O�S��#��D>^�e��<�kщ�L�bau��p��r� ��7���G�*mĩ�薙���!V��/, IO��,��Ӽ��^���b;MUka�%M2p��*���Y����j���3����:DOL�aI`�6�����R�0==����U��S /,��}p%Ќ8����9Q��IĎ��;/^ĭ=�|�:5is�(����D�b�ʄ�Q��Y��	|9����o���v�F>���},�X9"!e�>f�f�|��El�U���H��X>|�2*׮�_�twkk�_�¹g;;�˹B�ץ�B<_����� �<���m
�K9��8�O�����L'$RN�!��r�G��prJ��f�d��+�����O~���xOq�6�٬�n.,,���թ���E\X���h������~��/�9��MӤ}���bo���TgJ���W�&f�:�M�A���}�][]]Z\��L���'��V��}����YUJ%C���xCu������^�Sӳ���^�)l����yN��o���o��o��m�,+3	����SRj�ݐ�,��gb?�1r{�^��!��wbɓ"UD]���#�5�Z�d���ō�1r� ����}�թ>V=��:��N��yo�a�Q��"�����~s���=��G���ܸ�s}m��m�����a*�I�P6�h`�������v�v��/ο�.��/�5�&�]�C[���B�O�CL-�J>"9���Sٴ�8���t�<����ݙ�a/�t�l�{+k+f^;tt�V�����3nq��(�����e~����	?�n�!/�8Vt�1R�99���h2=99]�i���@¦r����,�~�����uh����b[�����>l��l�+e��	�Dx��i�j$�FA��(	}?�D�+�C��B�0�X�!��d D:�0�}����Jrx�P0�e�S���cQH��p ����ʌ��O?�ַ������
Ӌ�i��wF;�k��.Q�K�멊�m�-Uo�;w�>�����n����������H�O �4����d1��.�f��N�,����|�z�U�'ߔ��p�8m��cǎ5=����ޜ���q�?���&���f�+�&9�ŝY�3�p���)������ƣnE�E���e��쬲&:�P(��D:��t��;$Y��R�2��V�2Q�B���N�>q��1<7�j5Q�a`Ȟ����0� t��ۼ�������Y�)j���dܫN�}���{��4ggg���%<|#���F&�1�+���]R�g�Y��~�Ա�g��.V�w�����ƹs/�A�o����?���f���Z:vdqq����X���ԧ~�%�A�\����G>��s�k��_���������#��Љည�Z�j.b�>�l�w�W�]�o���G�8�j��nc�I�UV�^���R�(�ʪ�)$1'��1Z��; ���p�eJ�o�~$��$z��ٹ�v���/~q{{�*���bT�A<
@"z�\����p\(�[���� ����d�������0���~�(~��n���Q��#��$�^Y%j�030"�A�����l���>��t[�#7 �Ijר�L�w�h$^I,I^	 4*P-hgw�����W�� ��MC����}b�v��
�j�K��@B��zU�~ כ8���8.�=c}Z�vF��4kYb5��� b�T�85a����rmJ+
�N8mr���&+�1���y���m�p�MV���E�!�N�'[�.�~���H"���1DA$�$V'��H��Xua�uB�z�I+�������Rɫ�s�ݏN����]5�H��#A�8��2ak�9h���4q�E]1"NJ,5R)4T�X�D�F"wT�#�:B�3nVs�aE��V��M���!������OSߪ�:�t���@�?w��j�����R"߸��m��h�q�샱����u��Hdp�Ƴ�LȁJa�l��}��+g���S�ĕ+W�4��k���Ra�M����i�:� �#!_i$�h~Z�ܴ����y��:�:��E#�D���(��6�J��N��V������pub���Xfn��H�\`��~�bibf�5X����O�Q�����I��6sH��Lυ�[ԎA�/5��ı�����y�ƒA�kkFe~�8�C�D����K��n;_*��3!QBP��?F-l���K�I�ԉ3w�^�[���Ӿ��3���C?����p\m� ����Ӣ	�����&��1qS�R&	��	�)U�L$j�LE+�9D�0��kU<����R����y��oZQ��[M�px/��֍��Y�bJք5�S"ȳ&a���Y�rA/[Ƅ��ɉG�Ca↩d�i{vIB(� �j�V��n��XGÉ�M��arZ4Y�^S��x�"u;KE
mSv�P��ii:u�q�`Ύ��'��8	-bE�ޯ��v�Wg\@�tb������D���|���.��T����/�xҥD�%��KL���[��!!]�H�*�P����'z��ќlZN7c�#gSI�⮐)r�F51������3�Ӗ�`��(�����)Y9�	v"�x�Y75'�Ν;;@��A�(��RW���g��x���&UcL��9�ݝb>�����C���˗7�6���G���񤻾g�Sb���(K"Zd���ׯonnr���B�����2&Bm�B��W����x0�c�t��q��b�?>���]�^�g�"Bs�Ie
�|r6j�%�L���Ƹa!��(ײ#P��m���KS����La��zK��u�Pm��ĒYi��I���E �fL��pF�8n%3��	dħ��l6��S�2�+{�ZV͉0�Gh���t��'��p�A�6�3g��v���� �ۂ�Tt��z���ߑt�W~�W��gf���X.����n��������?�o���{'K���G~�w~?�9J:�V�������i߉��ޕ+�Ο?_�o����D�ʱ�nm� yp�}�(c�Y����Hp���:ʈS�x����W��I�+++���-� vxD�����|U��0?�$�,MEL�ڝ��5 �rm�PD?t"�ΛyU��{��ID�<���`Vn��f֡�r�0��"l+�R���F�Y��T$Ǎ���^3
�P��ҏ?t��v[T�ŗ�h7�\�3�,=�����s��A�C����1�#M�l����H*�/�-���*��h-�./���}��؇)�l|P��8*` ��6������4�Ni!RT"E��Y�� $e��^�����eŶ�a�� ����Qs��L�p_�%;5MHv�Zf4E,����
BCad�(�-���I|s����5>��MU��ۑE�L/�P,�]w����q*��9�cgƻ��T����t_TN�r�6��iEA*%3�E���|��7�g���.VȺ	��N$�h�`PH��$㩋C�8�a��B��(�J��Ⰼ���zW�\��KQ$��i�;�^�ŧT��hP��=A$�pr�6^$����lvF�LO"e��#ƾI"�0�c��U�PJx�c�ɭH"��A�K~��>^��	�p�<ϫ�&���g��z��ӧK�N������������]��|�8Y������j��[�$�/X�0T���:�u^rcM�B�4�����F�6Y5�K�z�qV;{;�j�n���j'�� ��{���7=3�[:�R;u�ęӲ��9S��x܎eY�y�*�1�%�a���?RqΓ���M¼(KJ�*�$��Y�M�#(^���IϞ(�'K�iHA??73�����:���B�TN�Wm{f~���C`��O5�8b0b��Un%�S�m�(�`J�Fy����R.��lSp֥��F(T]a�]Q���ӎa�`oj�(<��eW�GB_�sb4F���.A�-+�*9JC�!Z�3��Vb������W4�H���^��Q�=�.�Ȧt������������;S�d��˓��I�/�RO4�a*D��9%1*��6u�I�<��'��-N(*��c2�(��:G��0̜��*n ��c}�\�$�����B�4~������TP���S�N�#���|Ɉ5����7'�l�di�%���,��\8t�_���O��ݤ�'�.U�`���l���	��8n�^$�&+� FaC
���ڼI2����� �M%�W��d���.b��A񧸸���l(���N� ����6��G'�`�5��'�?������Pd<Ɂ/ì��h�����W-3��|��h��D<#qr���$WEv�K����~cQ�w��Q�
�`���!*�`�s��p�i��ūG]�������(֊cC��-ob��·�e��J珧�ﹿ����s�����,.-�vǙ�?{cm�����H�җ��*��_�o~�ێ9=Q�{�އ��NJ|N��Pl7��[������O>���ֆ���&���{^������58��0��U��u�Y�2��ey�7^?jp��������(�P��8A���A�K��0���S���Y;�qtif�*9�+*9j�Z;k,�F���w��vR��{�=
���"DR���#��CĈ��0fvJ�@�6W�y� �8"	�a��[v�"����5S#nlE�lC�M[�K�tZ��f��N������2�d�4�b��<n��7��#_�?
���,��{͖pr�N�#¹0���+j��J@'����*H�	�M�@IL�\�I�%d�x��g�f�D���6n�;�rz��0(L�>���\\4Ul�t#.�����*�H*%|�p�!ƔC��Hٙ	�
�l�]����h&n��<l	�n���]��/�`��jl�#:�J�@�#PD���������X�Dĩ|]�bGT'ڠIs��c	%±!�Hhbx�B��R�����k 9x��	�;�����+ yʨ���h��lIv�<��PR��4���XF���$�����ۊ#��15YE<7ǃh��PLY�pQ�Qxt����Р����$ ��z!�C�A)�-���}QDZhd��_���DzY�p�=Gm���BNJ�+�^��7�	g����n�۷�v�v���afi	K11Q-�s7�V66�s��f���^�8�s{sK�������NAH��V���]?�,��D�;��ӧ��/��R}k�ؑ#����+�Ӿ�;�C2��F��x[Z��L��Rt}f���� �ַ=����{�$��W&�٥�t���"6�7�ꮕu��K��o��B�}�Np�`�=��iH�^���
��İU�e��:AIҌBI�-'	Ub�3�|Ѷ
���i��*Y��t��m����OJ�&MN��v���ȋ��W
]٤Hs�T���{���/!�tm����S'
�EK�|��FL�B�F����uֈ8]<��"]E?˚��a	�M!b��2������y@/����z�x�I�f"����V�d�=/���f�1Q+---M�&.�|�����>xW�I��~�4�ϧT�K!��x~_S�.��@��s�"�ף4��r��H�Z���Nr�CR	��T\�yQ������F�.LO�(�	��G���E��F�0��������\YY9t�����nܸ1^`�o翊����	��3�iu�j)r�Z=z���#G���@L+Q�*�^3��h`mp:­h�b���� ��{aBm�������#����C����x/�>rk�i�����b{Ol9�b��d�Y))�V�$3Fֿ�S��Θ-���M(N��p
�)���������S����w;ϟo��EM1�3�L{ �T��q�sss�>	�	�HYLNQq/�򵂦fD(�}�$�-Ĭ�����QgD�Y��׊Y(Nϰ��b��/l�i�/|��o~�O��C��yY	��Πǭ�8<�bh�~���l�m?���~�,uj�X�Ƒ���?�������l����Z\\��1ucG���lo�ϝ�ҥ+_{�ɗ/�t��ʶ�y0�%>a%���͝�;o���7�\ϡ�
u�$w�P�.�!��������Q�?�
fd<�����Q�	c�H��f�GՋ�F��4��K��"�A�d�e�#o�n�E��l�2��^�G����'
֤�M�?�H%-����&�=&E�8>�VY�����z��54�`��K�@�'G#��b�LN���j����#M*�A��s1I����F8�j�F��" ���$� �4ĜQ�����x�R���~S��",��6t3�,���):���ǦH�I�E��ciB�R�1��q`Ө8���E4=,,)�?��
���=Պ�2q������I3�bߖ�G|,�	v����*Z�eN��� ���ML윀�Q�
�4�>I���,���0����}j��q
�U�WZ������oɦS�a��ʑ�"��6�9��z}q���0&�XR=մ�,*��C4mO�`iA@g x�t�$Dl�)��z������¯�Hs�-�UB9<jGT�)@�O8�'�;�d��[a�N<o��Hg����&� �
�1�����|��
���D�p{�[�T�,z�iG�;�{:.�J�*N�4F�&��VQڭ.1Jh�W�����}���%��o?FA��,jZ���$�M��u�|�T_{=� "�ۋK��춝�?������ \]]���8�յ�F{�q�xا�f܀�6�82�ئ���T���R�秣�i�v�����9 �r�a���Vw7����������Ŕ9A�P��έ�7-!�.��)MN ���hAL��#`P�TL܁��tO4�!c�U�"Q$�����ݦ�.{I�ȉe�I}���-��LWK�n��a�zZ�r�MD�Foukck���CsJ1/��x@���؎w7T��\aj��g����V����g�)���'�`LJ��)M%�B@-h�#�	 S�-�#vqo[���a��u���P�%�L��NߩoS�*��6�$����C�G/�������;�:iN/�:��(D��m�v=�P��km�����c��ɩ�׷���by��<� i��	��#�2�`�F)AkQ���N8���͋}�\�B�Z*��Y�8��l�=����P7����V+03?W�Q�2�#�ȈV��D�f����&�>��`S�~���.ˈt��<������VǏ����?������|�=��A+�l�)B��n��+LaI�x>ǬN�\�[[[���9y��iڢcVa6#b�)�(az�M'&D^z`,給)^u�\wd�	�3��q���4R��T��W
�fu���#�?�΍&���������m�,D������Q����e��>}��\� S%�1����#�����5W\ F����=��JE�mg��������}��~oo���h��l'^Z���:)��Г�	)E�^x������ƚa���++�ȯ*��;Iw��F��������g�s�I�z���Fs_�`��^/���r��o{�����G�mˀ�����9���Ϝ}�٧z��)U�n�����[|��o�خ��Z��76�$II;���֐��9��?c|(=���: �����x}�^�[[�n
�ɉh��E�I��U$
p���9�H�jJ��z�K�Q�ՁR�`�$-E�� [�[�L��8 ��	26�?T�o�4.G��Tj�4�R��7M�6�Id�1?2Ͳ�"�'>`|�J��QZ�iR@myD���7
9)I�x��O T�Q�.DN0��P�dCd�Ƒ)�6�p�	N�;��Rr�<J���S�B=�츀$��!R2�*RW�j;�?ǲmI*�|����H��#E��B=�u�aQT��G��
M�
s�o�<��Lp�T/�{��,UJ$na\d���i�mǁ�"a>=�@�	4���^L��W$����{)�cD��t��o*�4#�m5Q�!J�;���`#R��8��nj��=S�Qζ5�ur"o`���]�:K5��1�%�%��t�uȏ#���T�C���V�ޔ����b����0��l���� �(�?b��4���$*�#�)!����G�Y�(��+��D�ev�K����W���&�f��9�U���KZDÈ�ރ���mӢ$n��#��3&'+�~������] \;_\��x� vŤ�2�o �q	P%����z7}xm�5�N�#W��-��ǊB�'(�)~�:�@t�t�쳟��?�o�J��=��J�wqhx�xZ[����ff?���.�C�#�������#G���rs�����s����i��kvn��o܍Î�遳���B�n�E�0�4S�+����^�<���ZX*�J kq��׿��'��Q���@+8����s�9�ΟxK�!���������i�I�c/�9���p�,�h�$䉭L�"����ǞL�@D:} %@ڿ+���J����������Z�&�)�,������g�K���'�j4;��М��H�l�����ԝ�����ؤm��n�]��O�gf�P�cvJn�n��r�]&�UbwDD�9 �bJ�mMX��
��C*U��4��;�I�( j��r����%Up�+7K�R�MZ�M2�bF�H���8��jsX6^���uk�k�JJ�̇�N�w�v��]���ĥ���Mw������ڍխ�냹����r�0I����IL=���j�
�w����k35�V��n��縿Z��~�U~�!~�A2s$D�yx����]Ͱ��ݩ���o}���@Lo��6��QE���f�H;�]� 433�'�WR�g#1x9���QلJY���?��#ǎ~���aj.�fV9�g��&����I>=��7n���׾����衷�>��И�f��b�=7@{��3��[3�HF���3�_�g��R�e��m*~���D����{��Z���+ٗfU��8��JF��$��뮇�@��EM4�2=��Ў$��m�={��n�L��B*ߔ�[\Z�d��쬡���D�����̎��u�\���իI�dM����%:���P8D\�rĒ��8���H��f>t���g֐�9������~�0�����n79d�r�>`˕�W�\�.864q���4�_����?�����k�� �/	E;\K�������m��!����F�a��ǲ�Qooԟ�I4"�{!rg��X���J<�5d�~@�{jB��z���8"� ��P�!�N1�?`��-F�U��%*#��<�D'�8�}�8��=�4���Ee)�C /��nH؆�X$�U��$8��˚ФWb/ FdI�qJ}�8F�� KB(�C8CC㞈�9L#7�+�It�Єu&�Ŕ@���Ѐ0@ݾK������>����K�d_!0��V��JS0�` �+%?�PG
SŔMQ��9p�9	���bKq�,&RD)\�>�vB)��ǔ��"�g�Q�a�`�4p:F��Eu2��/q"D����k�[�y�0`�Wj?�xI����$�9U� �>LȔPx�#�ȕ.�*���9v�P�6v*��)����������5?F,��I���h�G:.�DҩOh;iA	_
��X��?�2����V<��T+Ib#Wd��x1�)	+i �Y'&��O�^S�Yg��*�&����N��i�C�íc��W,L��n��#�,iؼM%�\. �����4bϠ|*&�[�Di�n��t{b��U�+o�i��#'M����`������a'��	U�Dt>*��pe�C;;;++�:��]�ܟ/��!
U!��Dɯeʩ^to�=|�\ J��,�w#d����i���ٞ_^��K�����/�3�bQ�3�����ު����JE6ll��م�_���M�圢�{��C'��y3�(�����t�ؙ����S���՝V�y��[>�KN������k7V�,ckbr����T���l]�v��?��jp�"&P&!��&K�|�� ��O�a`a�H�Y��xnqsi��װ%5!#Bn�,bh�����R6�s�����+W��ח��k��q��Υ�!��U��b�Q�~��w})*�N�������������,�k��;��^�E�y�Y.OȰQ�D����K�����x2M�e�t8SGmQH��<j�r�A�݌e��R�i��'*jE�Wd�]�������̾x�P0�#�[�� ���ɷ��{z��I\C��Wby�VӁ�s�'N,=)�y5._�x����~�=���ݎ�u��1̦��Q[f��'r��3�{)�q&�2s�A��r����/�ڪ�ES,��̼Ѝ �+Y�`D�ŋ�~����҉��ܴ�j�x񥕕|5@T�I��
��,r�4v� $/��U,)�k6͒���a�~���6�ҥK��k������#�d,s|�L���>���.\�������+��"���W���u�p��a|ř3g�w�Ⅿ��wv�677qs�y晌ؚ#�������o���gZ��3b��Ƀ�2O@ƾ�%22����(e�k{\�U�p��$z���}�> �x������N�R��Uw���8y�-���|�F����G5];��R)��V}q`'����������>��A�l�6���컲I�ͳ2�3��P9dp0aC�z��خ3���ٖ��L�)�&�(�<w����n�
΃��k�m0r5���$�SP�� .n�i�z���M)��]S}�H���A�d�����F�n�jo ���0D�	
N�P?(��"b�
��}B�R�z�i$��!8��q��Cj��b-IE%"m��(������x�<3����F���'b�.��p?���-)uO�C m"�m��!#�~�l%��a�!W!+&'Čxd�C�����M,�(C[)�9<��s���H*U3���� nи�%e#���Ktʷ���"њNϩ�Lq��*Bpf�e���$#$5a�{4�tSU,��-m(��n���꩕�bϕXF�&���d�t��㐛E� 9;B��=Ӱgf&q���֠�z��:1�|A1tj��!��4���D�y��H*�K�טXqi,��;�Hh_R��6��o��4���6B�@׈��j4�ANN���6"�X&����aq���hl���.�z�D���Q��$:�S��G��X�4o>�i,�q�z1!����(%Ԕ��Se��b)N�Ur=�q�0�������hnGd�[�|���׀�O��|���¡�0�b��3��Wt��`�a5��g/�M�h�Չݖ3���mAϪr�rd��!�]*��|wwa6�X(����C,$6����&B�f���n�="�B����*��v�g�z�۝�AH������|�-��93=7;5{����bsw�.Oi��:�]0��ɳ/_�.�'�->������;w���E��o�(�Lת�|!��������O��_z������7/<w5?Y��m?���?��ϖ�3�@��������L�iʷ���`�]����/<�����N��ds����h��]�Գ�&�3�ЃO��9[�X;�xn(���M�H0�Q���h����{��s���C�aQ�,��SS�����4]���{��i EBJ��0�[Z��R<rT��tc������2l`�ԉ4��%���7w[V�LLNۓ�buR\L#SPD���74��������UDQ�	*��1	(��� *$D�B���~�K�����'�R��>}Pd0�vA�������r�J��X^u@�������ʦ���剩r8h���^��\8|DҬ��t��8�<ߝ�.t;�����?��gO?�Z�G<�f����T*^d4�{�b�4r^�j�r��(��y���뷁{gg+q\o6ھ�p�5ȩa����ٳg�������\qJR}E�bK���}�����p� @g�)'��qD�\ ��Pb$�j�����_XZ$ƹ�v���R ߣ�#��kkk7nܸ(^ <�M��'k��+\ڝwގ{�;��;O<�������ﾓa�ﻀg�<����U���� TC�ϊ���=PYM�i6g}tY��,5��!2;ڐC^n��Dr�3����Z�����2�\eZ����.�����/����s��m�>}��	�A|��
 �������>��35��˅C=���L���s��y�̉0�r|�������Ɓ́������bybj��Kd�֊u��B�܌c�0:�a�Yv���֩A[,��:_']��I�5�h��j��><�����k�K/�i��+��۪	�B�HX�0@�F�S�b�ˁ�S�:Q)*#1+�"�G
[D������Δ���
���q,�2>�9n=��H?��Zd��=N�.!{'��T��J�81uCF��
��h�KF��xn�Q8�QSb��Vu@� ���*������p|J>��E�h�E�äf�5��B$@-�~�*�{{r�Ǣ"k�E�ʬ�t�a���������o*�V�\� �D�!�)�I�0Ӹ��D��g2	���EnD:2"'Q�[����	�"�$+������'̢��=�O�Ē�Ps����s@G�?�5bӍjIRĮj��C�q:Q���{X�!�t&���Z��i�_r).��rN�t���=�q�d�}7j���)-Wj�nz�Q&TG(K���e����>��|y��i-'�p���T2}�����ng;!�S�Ҹ�/�8�iK�-2U��i�����͌!)�����, @�B6-�LI*�X%ͥ��>N�.���ۦf$�܏�b����S�/Wҍ���@)l�kST�dG�27t�1nb��p�@�a�z���f�R=����M��2M�a��;��&ن�If��T�!��j�]F:���lq9�	�Q�b���;��,�;���B�N�vc�턽P�.hn}��酉I����󢨛�z�Y1
��&�/�d3N5���ƖBQ�T�V.I�@L�A��R�0�}!���
B�CH�h���;N�n����Rp˻$�s3��'��^1_Aȫ"*-����?���{+ʪ��|��(_�t�O�%�*������j�����_�l�ؑ;��p�ݐ(�>Wеj$��߁*MK�YA��������Z�W�����;���1�ӾQ�:������/K�f9��V��{��O=�-b@�~B��Hя��Qr)�c*���
�n����K�{�O��'�41I�VN&K��ٙ�[W�A gë�XF�	�ֈbb�P��%��N��¡�#5x��.!�<<����q��
���<Ů,�=/)i�h V��z⪩t���ɣ:1���]̘�93�P��9�L�&Ǌ���~��4�S���M#w*�Mc9Gti�����2U�D����U�ҐTzbQ�d����#8dUr�p�\���I���NNO�9��& �,"���������n��{�<�i��[������c��,P�0@6���[��f^G4��`��*���eX~0i���܉�Rq��6U�!-+�ln�;����yә��-ې�.����s��L(�?thaq��/�������<͈vw6f&g�
¹�~8=5�s�%yo�'�����ǎZ�����ۈzSo����������9s9u�Lo���6�j�R��?�����w�}VՈ�G��0|K��U�`4�����O`g�o��1�b7NV&������3�;v�taZ��?���_��ׯ^�ʊ�,!��|���>s�5�DL��z���N��h���8%�k��l|V��Y�&�'�kaG�*Y��@��kA,�C��#�ь���xW0��"��^������d��X�S7b������ɣGy�����}��o�������ovv6�+|�O}���\X��8��\�|���{׻ޅͰ��4�l���r�����_���O}*#����lN���ʲ:Xւ��h�7���^	69�AՔ�CRiʚ8Q��cs!��a��Q��P3�)���y�5��@��0s�tFK(�O���W�p�*+��D:)��Q�Fr��іRo�"&�.6Z'�0J\"ST&4"W�����"')��";@|��e�&����J�M�N������?56�fҤב�N�ƴ�x�H�&�["�?cyDJf�T5��K�Eitz�����L�T��)cD���R���� 2�}'���,3G}â?M�[�w��&4|��h���s�R���w���v��-V��o:V�&�D�Fg��FsX�{f�T�Y�z͍�����`(���HҔ,�t��U�����r��M����9����N��I�,�=<Y.��j��w<��ޞ�+���iD�a:n�=���"��9�Z�f����z
Vtי����k55Y�i��t���rn��N����
^��U��˓QJޠUo�o��ۨ�|��`�u�@StiHN�Y�yhi�Ȓa��!���zc��1�֬��C��9n���� ��[�dy��
}����"��`�Ҽ�`�Qe%K"�7�RZ��1.�7Y�n����L��mo���m���ܱ�K�J1�T�F�v���7ֺ�v�dLN����؉���F��PyGH"���o'@*��92y��bA&Oy��n�վ}ɼ�Ӈ��w�~}����v�W_�2M���?���)^��uI�ߧ�(:>������\5������l�p5>yt&���K�˻�����5�4&�6b���~��\�;y���n�k����w����s��ڥ|aS���Y
7�����"j��#c�i���[���I�q�*�tZm�.C�c��iߘ�Q���)s%�F���Q2�v!�k�K��3����^��wN�:1U��#�l�+��	��ǳ|\���+���F�7.^�����>���
��j���cv��u���|�$}�T��-�p�]Y�T���*Q�꺱�� |�f|b���܃>�c?�c�2��b]c���癗�ٖ�)J�s2���G��/�T�ŀ�h��R�������
��'1Y�5�|2��� �ŢR(�tɒ���kd�yb�S�8��T�b��mլ*R�($4Mw�w�8�c
(�τ�-�G�#�E*�N�q���,����<�� xnnnc}��45%+�/F�|��E��+++���][\�����Ur+��ȧ�b]�iJ�N��w_>~��du
���ʹ
)��%��Y� �M��{�I&8m,Z�q� `��t4])揾��_|��_y�˅"|S�9�0�uw�Z�~���)a�V~�[���w>&���'#�'T��)؂���OO��$.�&�V��+�����������>}�ɯ�#�e���>����S����_��_mll9r{�;v)��o��T�� /���]�����`I�V*�p�Wy(`rff�?�_�.Sca����eMn�8�� I�axwe�5c��k�ՠe6�@�ݫ8�M���N9I���b	�LL�>}K�-���}�Ś���X+��G��#^
EY]]�#������o�;������8�o;|�p�Z�3���&r{%a�4F�8j̡I�l�W��S�+%R�D
������cQn�S����&��'9#��n%����6��a�"�·%>�Ds�h�OP��X�"�i#�.l*S�r~@��џs����Pp<Q��k��b	j�$� �B<�����6T�SԶ�a�*d?@��:`� B?B��VTa�T�~���i���N|�C���~zcs{֛���c�k��U)���m�sSg�{���7^Z8���Z�o�Ϝ�re�+�Y{�a�q���LXX5����ܣ����{(���L��T���:���I�@�9S�DR��e��������>�����뱽^{F�wtd[HK")1� I����F��Օ���o�C�AR$W�h�a��Ө~U���������W=|li�V�����{�曯�ۤÅӳ�}��T�:?{�𑗞:�8LaC�$�3/��k�X`Cjav=���~�� ��4���گ�_��g�x|||i�`�k�����]�$��4������3O�|�šbٌ�����4���/L6��&���-q<��$p�mO��\5	���1���7�S�]�#�=3t�|�Sܲ����8�9�H��
+�%3/�8s�ȫ�%WHt�a����(��������0:�/���EAW��T�������y��Щs�����o�=��M�����p�f����_>t�q��l>VX���/�=�«��ˈX�����)�.�آ��r0�w޾�s�zoya�yԮp����޿w���uf�K�T<�R󱎳gN:�ӡӧe1\�~},�o�w~�|����+ؑ�E�I��JQj`��?x�]��Ώ�{��U��-[�����E�O�T��u=H�
��ڡ�y�*���DgO �S3��?rίq�A�9�-'e[k�K�6r���X�������#�������޸�}7�Y�9���ͺ���'>�B�X�8{׶5s�\ߪ�Ξ���щE%��vx�����=eE�����i��M[L�{�v�t�Αp� I�ja)�<��&�<>ڎ��b��-.˥���������E�k�,M�,N+���f��]�6P���?��4 lÞ�a*���`a)h�����n�D���ٹ����d:�qsJ	���eE���k�����=����b��@�,�?#�e���6"��5$5���U�G6)����GG2[1}] 	S������P������x�2 ��ȺlXE�NTD�OM �Z�fx�G��=	q	�
�X1�bЉ !&9�McCJoЫ7oQx���.� �o��εz���/�4�l@�2m�]�8�<���	 ���������a ��">"��2�]2L��[��z��-;v1Ɍmz��ך�#�H�E�՘J�Y^N�2�&Y���D���2ف��o��{o�Uurb�'�{��3�Q��y�a���f0xhI�&*qIEGBj�m�:,rA�	�C� T7@�i4'nٺ��[n<r�����fn��{����&��H�8�x:'i�T*Eot�����s��@9 ����*<D*� p��_ ��(
M���ܲfϲs��o\��Er�5�(}�Yo'	Q�,�?��;��E������
F��;z�W���/�Q����ȋ�_����RT9F�?Xt|���O>��sϭ]��P(��`3/\� �f#GP� �N���%�C��F�w��	�@&ꥡqU&д�i4a'N�Q��x	9��r]p��T�s��b	��'��R�o�q�"i�1pa���|�������PUL�"y@I�Ds�Ĺ`�����H�Ve&jO�Y��aa�2M[�d<A�(٦nX��i���ô��j������e	7�u!�{��Q)s��,|��a[z�H%���?���Ǟyl�c��~�W\�?ӑ^�.O��.4:2Z�w������|Oq���W^?3�9��t��b���AK�O!5��0}tyM������o�q����#/����0�����5��>w���-ړ�k6��w��{vߴi�M����|��=��R����y��xE��>��fD��g� 0��bz����p�-�}�������\��O}v��KK�c/=��qN���۰a`��7��z���Z�9��r�ħU	��|��Ai7��b|�ॵd|Fݾ{�u7��9�����Ś�+����� �KG_;pʬ�*�ؿq�{n����S�����K��սkbRB�c�"�f�EҢ��(��`��i7�I"ծ�k�l��w2<1��O��}~���щ�N�
�f�+=]���sͧ��	���G�9�ҙ�۽Z���YE���rJ��(6����0�s!�p��n���+o��O���^==��O~�O��`��xq���L,����ܵy�UW�꺫���#?����7gR�|"���r,lájs��zIذX0���ۮ���\Z����Sw������]����}�k��x���T�p��w=��;�ܰw��W}���^�M�����ߕ�Y";J|�Dӂ�4��*g��xݺu[�l:5:9ۙ��w�m��xkG��s���P-g���>�w��۾���N9�H����7��w�:Yn�iؼ :$�浰�#|: ���,q(b�+��%(7��o�W�S�h�>*��<�T���"�����8</�6��}����'GΝ�x�����=��ށ-��׭��^��:��S��Â��.l(b��$�@�m�Og3�eV��zÊe��lڞ��eU�o�\��-���g;2�,kԍ���5�]��R�3�Uk7`Ѐ!��h06_
i��Ft��[�RV.G���Y�^F����@���Kr�$�cs����QdF�o�|ȑ�a�g7"p�b�q+εt��y�wM��X^E�)��X.P%QN0��XX&=�6�]�$��4��!�Qt�óX���!`e�b֥���/�w��+�ڙ����p��2�f��d'x�R!q��v%��h�h�J �N&�###����2��,��bE����J+�p���P��(q��̋ a:*����W�Pƚ�q �u�����޵��w^��=, :9s��'�����3�� �Vk��a��ǈX��2AXA��11�E�)�"�2��D�'R|0�`����������x�b;��<��n��$DEQ��*�=Q�ɬ�,8���)���Q�I�B�L�
L{d d���f�w�	���/�OQ���@]�� �2�;��QL���a{��/z�QG�HJ.2D+KtX��v9�Y!����;E](WD��h0
8$�8��]�����'�D��7Ce����G}}}�6m��D������� %�Q'%�mt��A�P�>������.*�Ge͗G�%���y��J�:��=���6�0 i�t�4\NQ2�t.�{P-WR��alׂi����Z��_L�;���^�$�.�ѵQtY�\C�0)_��YL?N��i�`�{X�Lzy�����<�כQM�LM��s떞��T&W7�j�aX���8`�����I�y�����h]���Ex�P��m��,W�\[5�_*/��ҡ����}7�z�m����?������Ό��1����ᦽ����;nݾC̲;���Zru'pt2�xm�Gt�\���爬��k�r��Ń:�t����s�MO8�|��.��U��H��������}���|���x�,?�䣦e�(��-�ɠ��H
�v5��E|8P��@Me���L����+n���=���������"\xWߚd��[��o��w������g�{�R.':���4`&Tl�$?p��c�5Z>��aA���Tݶ���C�?w�}��C�������������Y�������?s���q��4=屇ؘ�d�ݕ��ʇ[����u�������KrmYLds��S�9�~��;���b]������yrb�f�
O�sW]���_���nIv������\^����װ�I���Ն��kHU��++�m�711�ܱ�=�?��;^���_����#����&q=ݩ>t�o��'����|���CS��W����?�@ھ������*ՐIg<�Ӄϟ�������~����×�����C�g9v��Cg?x������[������Ɔ�v�I�K�"&�cGUz>�Ţ�@^#>@50ހ6f&�^=q�����Gn��cg���_:p��RIWd~��uw�u띷���_VT�̱��r<[�)��cE5�h:�w6ҡ;5]��4��A\�"%3��$D����{��Ŏ�xE}���b��(�p��w&@m>Ɨ%�+�WO��p�8=56t&_H~�C�t�W��Q$�3j㩤�g׭�XO�a[��v^��n]7O������B}���6���5A! �<?5��=q����|!��2�;j��Z�^�g��Dg>-˰��Y��J�{��د���|�Q���_&�Ѳ�?��)d�1㝶����+,�sE	(��6Pcq9�.��Ȗ���T���c|�W4�E�n����&
~�c������v�ׁS���<�p��J��cX�9��L����4�.A�������t��a��g<iW@�-W��� �Fæ`ڸ��h�a�T�i�4Y�}�������v���[(`�T*�Oo����!�	��NH(.,��g�[�kc����\1�$�]�̈�Z,�s��(��L/��$��5}F-����F-�TG���>kc���������8}��-�ޙJ0?�j��������Bg�����jʲS� �e�Y@r0gdE���$; ̜���A�gF��:���`��)�>O�>��\hff<j��ϋ�5����tuua�e]���T�و��J���o�1 ��b�J���_ɹ<i�usO��<Vdܽ�uG,Y�߉�ĊYW.��i��e�;��߸q#�$�:��eA�[/��7�"�����0ڔ�F:���]�����qzj���Zpm4۞�M�V�N:Ydz{n��ֻ�^����L���������D5�rP� lj�#�(�cG�,�غ��o�CAQM*�D,��AI2��D�okH]&!�A^�dbj�A�M\+:�p�Tf��^�399y����\��`㶭Z2���||lr��]?��w��S��R���E��*z7��{��h`�墢�dqҵښu�^(.�8Q���ؽ�ʛo��셱���<���m"R��tK_b|qzv�ĉ�^����n����X�̗5��M�o%�a�3��P�������ј��.��럸�����G�������D:&�LBV��3rz���JN=�������U���x�/c�{���0�k�/���&\��&$Q�7*�Ϝ����}|�����W���~���JR�c2�!eaz��菎M��Ɵ~����}~|���(�B��>�VI���Ԍ��{���eA�^�:qˍ{?�{�7rq�w?�G��;hz(Ju�b.����?=z�ſ��߿�ԧ�O<�c�9ޗd���״�h�R��L�	x�< B�cZ�rim_ׯ��KK���|�_=`&"�/;��L���<w@7��㣿��7�滰���Se�E��dZ�о-ї,( Lɇͩ:99�f���_���ϗ���}0GR��1����Ȍ���WK����v�>R�U�Ǖ8IEǤF�KǪ��H�+��[;%�흚�����7��������������D�` C��ٙů~u�������m�����g��t*���5O���ē�%�b�n���$EL���%H��׫ �?����r�/�౧�������.ʉ��t����=������~������g'ύ��d�T���ɚ���^㸴������]���;�rD����=�,�L4ǌYn�'r, ( �	-���زy�c�H6��uA��/�>���훺>62rյ޵go,S0�c+��՛�
c�b�����
�45�/����Y�Rq%�E'����$W5����,H��I�W���ŗ��ݳ�6��f�V.bKD��S������S��'���� �t�7�_@����L���t||ꩧ�lX���i�8PoK}9����J���<jI:��8(��H< I�Q*��l��5��]5�%Ҿ��(�)��YXsǠT'�S��iJ���\ ���]�GqƐ�S���{x��Ψ����V��-��Wh��^qT�h��N=���t8��NZ7�a��u�S0��7u����~��>	0e~~~nn��F��'�?	�ak�NT�O�z��G~8W4�P�_,ի����"���q��}�L��nO=s�[�|�2����Woذ.2��^:����ӵfs*�q���W��;/~���Inh����0����nd~~����#�v����ݵu��D"�9v�Շ���_��������������S���厘�ƾE\���8`���-=,������'�����4 7K낢�LY
m�N���Rt�o5$ )R�o�^���\ϡO߈
���@ӊ1l�$�R
����"y�.I �gggW�Z�����Q.Ǵ���J��P���H�F	>K���(;���;�u����_�(ҙhe�!g�G@�)	���;vl}���������5M����S�ZU��'������l�K���b!plF7��k�VI�x	��F��[�[��5=xQ����N�-ݤG*���u��⚦(��T:�D�l����*�{p�ƅӴ��oKK�\GGgAV�T&����O72�����g�B�5T�bA���Y���4)n9�)LNN�����}}=�r�+����Oî�i
��'b�P�7���?�_��k����;3[v�9?"2��!��/�~�V��z�ЌTʚD�F�:�����;�������� �d�^ץ��G�#ȍ��׿�X.���?���o��@�,;���`�!�_Q)�cWHU.�1�|OP�����g��kv�~�{�������vۍ�`%7�%VXU^�}�+�\�i��>~Ŏ���|뇓ï�`��{Ԏc*#��^�~jlA���t���(���w���֗��/>�,X�-f8�z���l��kS�~������ot��M��p�Z2ƺXɈ׮s�ZQWƣ��@9A�r�ѩw�q뺵����ﻡ�%⮭+�$lخ-LU��m^ݻ}�c�/k�߮7�M�b��H��4b�qO$�X@vV�R펛o���}��=��SU�4��ǒj2��T������k�_s���W�,���x�%�/9@�~��]��}��Pع��U���o?��/}��f�b"�Ħ�׊	r�7�4�ǟ?�w�����w��_�����,�K(�C�?T �?���H��R!M͟����ƛ��x�������٥l6�lX��%cZ�i���}�����'>�������C�ne������*�2�\$B	�}��'ȶv)�%3Ek��	0ǄoȢ��^���Hߠ�~�0܋(�۶m۴e�n<���G_|~d�B.����Z*Ws�-�5�`��K,/JB<�p�E�f�+�\�ö�lLKچ�8���bū�n����1���ёΤ�[����>4=;ӷ0�N&�\"��	�j������-[�uX+3�B���R;��;Ie{��8�^"���}�嗏=��O}�������	��r� �j= u�����W��/�kKS��y�&֑X5 ���r���Ten��l�����!���@��,].�͈����[8��c�l�Z���8A��]i,��=�)���0�>T�'��&+��q�gsB+1	B���(1	��>�%�E��:y�q퉼��xʂ��+ � �M������-�/�·b�h�B���Qup���ɹ��w~��a�����?;�cp��^T���Ӵk��O<���?b6�x\�x�UO<�� ({h����_x��W3��������5I�|����w���'kտ��z��  �l�ś�[�����k�y���e<O�SK��d2�ٙ�������MV��6+����R�Jߧ9H�a��O:��'%H���ˣ�}�tzЇN�5�ZQ�����������B��
�5��U���<+�L�k��]ξV$ ����#=:�M��0�h2pGG�Eu��A��(K7P�v�]D�-�#E#��yD�>_��ʍ��z��â�c�MI�Lא幐@��T2��~���3K��891/���|>۝)8�566r��W&��\�H;1-�R\Mr�lqa��蘂]S�(Q�U�c���]-�^-��v��V�D2Wi��$	�|y"�Z���#�܂���a�]�~PM$����>$��=��#�����(�M�z�$��[���$��j����/j�eE^/C�]�˦*�����W&���: ,�~��l���X�=ؕ���6f�]���;��Ӈ6��.t��J��q[7��ö?~�&���;e�.��a�a�3���s�g[_�߿���3�D����z�B�]X���i��O�uv��]�D��T�1��$Nx����3�
� �D�����
X9�I�\�J��Ǿ���B-��U�;�#�,5*���g3ɾJu��?��u�
[��v�˖P��`AG�R.XH˶��*ڥ��n��W�P�����������{2�ʞ��ئ���'�i�0W�F��:x��w�ݹ�����'9x�t��O�=>�]r��^R.֬�:;�W�~�����PNO� x��N�Vɼ��ɓ�O=yx���W��g�ؾ���'�5�s�M�(*��ݓM�g �c5&��ba ��U��s?}�?��R�!h
C��&�CT��zs��3c3}�W�ܶkwiv�޴)�[�6P���a�K|���{﻿<[�ۯ|��sS��4<U����Wk{w]1�q��#���S��]�����w2?��i��?��[��[��ZM������k7�:�N]���%��\>m4���
.IwB��eӥJ������}Ǧ�������n�b1ն̈́��4�i�I�Q{<�$�4F����������0��  �`� ����<�"��x<	� @�Y*Wҩ$��`!+�/?~�� �7=;�Le�{{PDM�ӹ�^m���LN��;'ذ^�f:b��ؔ���_,,C�w����m�M$�� 2�_��r8>��V�%|F\XjL����'�R[c�\����x�5_��/>u���촪�aO$pD$���������)���Gݺ(1oK4�:�s�"��-�d����j�j&XNmrf����Q�%��kֈJGw^�ư+s�C���1Z��VX���뵱������ݜ��$��� �3'Oc9i͚�0�|�dxl$��Q@�I�'	 �o�6��)<�A^��<�bk`�ZV�	�n������I���@Z+��"��s�͇Ѡ�8˒'Hԋ�"�ڨ��;�b,�U)D�$}�
'k�LB-��#�3��	GU1M%���S��ow��}pK�rS�#"����M}���%]��.�X�ߙ�bA�U���y�,�_`;0�4U'�<h=�P�|x�����������tu����Cf��%A��xnn����� Y�&�i�)"�zs���-�j/��CM�Btۍ���%j�-�����(���VQzCA'iV�2˺s�y�/4��~zAX�������E�U���#��]-Ro��{-������aS�N;�� FR��f~�Ô&R6�,��QzC��-���)
��϶W��;�HХD�=6�%'���B�UJ�d˳I(2l!�6�ر3��mZܙs�����56o�]�z�����f?{����r���t��C
�Z8Q___����J�d���-��k}���n[0\�$�p���eƠ4\9���-�(E1.b"Չ8[ +R.JM�����;w�s����n�@��^S�֯_�����a0�:��5"�>��h�{���Ei,^�����n#+s<K�J8��}}�l9v��Ӈ��2v-�_[�{! ���V�f�г��mga}��}�1t���� �a`�cI�Ґ��PGp9ˡ;40)����6��\���ΜVX�lT��8v�T,�"'xu�[��p������wo�X?i�(��{u!�m΢��UI���G�H��>L9a�BV4��'�;�p��`�l+h���f�Pe���Ǉ�O��o���m[vn<���K�Y��eUl;���2	�	����Z���=X�T.6�f�#{���<��\�$��rR�\{mW^�.#�<v�?=:�p��^�r{ז��2�{x.&Y�j���#�Ֆm�5��ka�?�On�%zjg|������'�}qn���Bӳ<x�"o^*�a]g~~�W|��9162���7y/�H�����b��!Ĵg�F�_�{����4,���{�S�������R4���o���QKǅ��N0Xa0�����ty�ւa���Vva1�E)�hZ�93��u��n���`\ܠ3���������q�6����M�[e7��)m�W��裧.��:�S�^��9%�7m8L;��"�[yq����'���-z! T�m�n4��<�ݣg�BIY*5$>����Yj,ńq&�kM��Oܼ��log�V����:�ٰM� �CY��������.��=* ���bV%&�<I��Y��\/4Ikc��U�%a�:��K�Q��U��,�j%�Sp�߿N
PUB���b!���n����l����g��D��5����Bs��k;�E�E��9���츢��VMM�f����V6_����T�LNey;�����j�c���$��%T�����W�9~������]{=?�h� i{&si2�'�l}�3W�t��6����
���tu���8]��à�z��#aSX�'(�pL��K)�=s�44�c렠�CgF�N���2]幥�����ܖ�븀�x~��B)c�-[���F��ܖ�]@��'��|�7#���[�u�
������?����T���ʇ��i��	`011l�.f�0^<��՝L����X�r�p>0�&��f=0M��Y Q����Dtu��e��tvbf��۪�pp��׎A)���D"c��H�������u8[���8���b\�w
QS�Wb	�g�JUd����J�F��C��y�g/~�a���e�)k�����D����D�ERb�Y��@�YoX��=���D�t�MB%YUb1lY��֍�ϿI�!I�tl�r�1���I�ɵ�0�Xt�D�B��)O{��[�|/��1T��P�I"	q�l�tV4!�;��];�h��a�KK�MIVׇ���e����9Q{꒏"� DED턤����s��0�ak�S$��I�����5\t�E)dQ2[�!)|�/۴�?J�-�H\ZD����c�&���D8z����	CE�����V0Jx�����L9ѶݷHw۳�i6��Р
�1Y����f;��xgnv�Dߊ�6z�*����7ݍ}����b� 8����z��/<�G��f��.Xl�y�+�&g��WUe���I����@�3�2|?�٦	;��[Sr�:���x�+��J����
>Ӛ�����q�|>.���@~l�e���9b8�s�7�J6;c`�$�4ZU��}ݷ�~���*��Q-��J�5P�ț ��<}��G5�F,��isX��dai@p�}⺤�l�>�>���w�QK��������)���K5<��\�5�W���W��J<�(
&y� &ZF�W̷Y�3�MO���X^�Q�Hu���yOy9c@S�H���dJ|�ݡ���/Lt616�V�BXC�g�f�3� ���R ��� �8�m*������Z��1R��چ�lBR񔢊�_|��ON��]C�tLT��1�q"��ؓ<?.b{�.A�0R��3 �C]Ȑ�/eX�����$l��8;r��ɥ҂��Л��ӱ3��x��	 d��k�̩�|_ZM�M�^�<��&���sq���һ
p W�}Y*������S�O׫�"�|�Bѳ��Ó,+�Uj������B\Q��-5m��l1|�g�Y�0��cLNN�]M��;����UM���ް2i��+滕�`{�"g&��<=1�m`�0�SC�篘>m/�� �&�r�|���sEIM�Vo�}.�{-#/6f_<a=}\M��R�i�`���4��E�Z�������HCx�:�q�%��}:��]<wff�4܃ȅ��z�p_p�IU��Z�7�˰i5��Ӳ�%��D"��`���;.VX����vV�:-JH�0�F���[^��m��D6r�S��N/�(v�`��19=mZ&l�NÎ'���g����xvU�QD�&�P�C�|�HFr��y��%X ��?��`2K�İ<9MV$�1{zz4E�4�P�)����Ţ�i0@�z	Vz&�s�칉���0�ka��L���XӰl��`�m4�4�cH�0���ֳ���;� �
r`B�8$���|hY ��ގ�5���a��K���{�l��8=��^a�:�K�nq~>lVY�
3��X"��_��co��~�/�'B�B��p�,�4&�������_�^.�� <wӕ;WlC
 ���d^y@����x��*yD�����s�l(�6?!�T���0��X"��Z�.K�彽:�v�/Z���yA�X�GZ�p��9���f\���!Q8ۘ`�c�F������av�`e���}�v$�XׁI��c�7�1G�Qb�z�v�X\`Lb�+�c��:�r`���j���c�Z�`���$��f��`BYR	�w�5�cڞ���i5��!c!�Z�_W��4<�Y�����1����fi���`][�����K�a�SvAW�JGrp�x���xȊ$"BY��C#6ʌ8L��W� E>�˷��CQ|�y�>�p,'�by'f���&��/�,��v�X,N�:$A�v��LX�O�0\7�BF0����� ���J�(�}<�xA�o`�J�
RP�� tժ�].�Y���כ��2�b'�Hm߾}��������ˇ\:��4����(��\.+�B@Sc@<L��e;R�4��PX��	{4g63iZm�����b�5Pzl��x8�1�RqqQd8*��7��5���^*���&��pc%�ª-�c���Q�'�)�o�<ƚlT���;�	L�v;��d�������W��MX�d~���O��cZJK���K�v�ޒ�{WS���#�?��"'�m��4��)ʞ�\ºj�UV/Wj�
O`��
��z ��}lB(�]Kw����Iв'��ByZ���6�,�$�L�h��� :%60��V�1Mk��+~`��T%ɲp\�P��'{��NҰω����b�~�F
C�h�xV��,�O���³1B(�c$^z'z�a��l�h,yM�.�����%0�{1��,��J�;Ұd���Ҹ@�.�'�kC�E��ۅ-�^�x�%֫U�N��El�a�u׬�!���J"'�pPQD
�S���:]z�@�XǷ�q���0`�,3p<K��ᙂ��]i����@R�J�	`���#$��2Չ�݈p[$�\�L]�^��r�� T�,�8z�e?���� V�$d����uuj\yf��(�.&���)��M��r����\^�'������e`;v=;�V��2p��j�eӀ=Щ荪�ç�.WD��ig�eƎt(�$,`��8K1:�Jɱ���l�KMoq�7�Ԫ����%��J��55�w���V`�y����L��a- ���h����6z'��(�^0�'�]�fiˉ(o.���:�Q<DT�$��L�f�$P����-�='&Y���nz�R�EQP%�x�C��\Ӭ"��� I�b9PVZ�KT`_"~k��H�$����B�!���w��^3�f�@qq�@�s��P�J2�mOc�����#���n��6�ζ.�y�O%b��%"�F9&��	�Q�d�&k� $b>�U�WzH#KT� ��J���[���t1�����̱�L�7]}A�g��.&L�b�X:�el�Q��q�g#�x�Vrk|6�q
㳀���'2J�V�Z�Z�5t^�$˨�ny���ܱ���� �`�I�\A�i�м6lI�O��3�T"Q�4pn��$R��xI�\@6X��bq~q�C��w�_D\��Ǽ	r}�ø��芥���M}
��Ӳ���J�s�u]ö0� l��̦ך�dԘV��*K%�T9�/ɀ� �U%�XםTLN&�4E�P(H�P.U¡AFI	��n�<��SX�v]<�{a�2�͉ɱ����#י�w���\,���Z2��]��a���b���#b��j;2�\�il�l��+�E☮�n"�e�T)�����PҭT*'N���jQ�P#�5Fj�4@E��7��
@�1�(kn�`��'ۑ��T\��}9��˩��B��'�m[QD�W{��%Ǣ�%10�@II%��XF��0�ӘMJ�Q����Ƶj�#�^Y��b0�l+,�*P`����k��l�j��v���bA�I�P�}<<#�Ա\�5ȃS�FH��$ՋDX}�� �`zi�0L�������<�u�R�l�F�\]�nQ��ǫTj4M.�3s�J��%� ��S<՘��t�bhPf0p���0x�\.�،_�����aaRL�9�0	����Q����v%U���z�jqQ��nB�;��01�xad���'�ya=��"F�˽�hU-��Hș�no�t.I��;D����]$B�Wj�6b�.dc���+���l&�Be��!�a���m��n�AŦ޼jǾ�d�Z����⎑9�f�M�k��(�A�GCȞ�$@�����TL\4���3o������+C�­���ܶ�����P\E֩��8�ؗ�h����(Y.z�YN�LP��5�'&Ó��0l��Ť��՞Scj"��T�j��=���.�>��[��ڠKM.���~P8$���A}8��$�L�/�f(KJ,��lif�4�K���⮭Y;=7�X��bJ�B���X�~��)q�a�B��ֳ�b^�d���­�{ ����;�x��6�i�y��b}bvf`U��7v�����%S�s��7���Q�H�2ū�\�+�,�f}C�	�k"l�l*�s�*|��=�n�|��GGW��8���6B<�ؐ�x���I8�Q�I��=�\��Ϟc%��l�*�����\Fs*��.ӑ�l\[oTa`�̪O&R��2-oE*#�!B���m�,�%E���H�_��� '�g�d���fe��k̪��j�R��5��t|ff N�X�-_�c��ʊ��v��Ʊ4@��/û$��,
i��#�y�Y�I�ʄo�>!X.����4�nE4�	�Ӂח�-QW{�6�kF�)�r\ęrM�8��@�S�Sa}�Nm[�ҁ�8���N��H�d�x�-y4+���	jk
 ����x����aT8�m��,�=�]���Y��+P��rh��	(,����R�L_1L�I"�bL%�[�T	L��[��a[u�D�����≁�&6oU��cRl¥�Iĵ�l����SgC7nW�~�6�&�5
1�+i��ا]oz�%�
}N��u�vi��;�M�vw���0�w|!P2�W�qM�2lVc���\&�`����[hR1h�ێ����W�N���ۛ�ǒ�Z�p���e�vCoR����8��Q�ܛ��l�R�J�:��u����P^n�x*�e��F1��9����U vrL+W+�z�(��,ۅ��`�``U/��f�� ������K���Y��L&E�Z��6X��ۻj��M�dC@��hV��'&��:�O0�dY���9???���$�t���/8��O?K�R�
�@1g����߿?���1��j.�??11��󝞞>�[Lӌ����մ8��%#�L�(���rMݜ���+�V���F�'�"3�K�*�E~�����D��"�$ʸk��� �h�{��K�f9�9+#]��m���VKO�~��K��D�2�����#�օgc�'	7h����Q ��	.����T`sH|�8�솞�G���['y�:h��_�Vŵ�ؓ�j���9���ӳ���<\�B��7,�G8Owa��&=�i��gΟq-��� �GҺ����z.��Ҵ���U`��M��k&)j,M����ӆ�4X�fZ��'�"`9���X���<iT����pR���ۊ�c���Vttz�n�1�i�1���dϊe��&�-��4�X'�}/�e�u���I��QP�U�E�fڻ��T�e?wٻ�^�vhEǴHy,
�n���uO��S�eWO�`�Cs��C�y��(�i���a�]MO�?���tj�ȴg�ea��d�@nhl���#.�J�������1j�#])(U�Q5�D�	O�u�e�xܲpr�,�fw>}��oY�:{�<�-� cZj�1^��ԺM�cO0"V��a&�-�:&q�@*��z�b�V�a;U'�� �b2��8�Q��|��5��|���JqU_���pHg5��H�Xj�W�[�vXQ508�Wz{*��:.�$z�1)�^"U�fe��vm�m7]_*�O�j_!H�0ML�o!�66���s��fE�jp����~�T'�P�,.%�aئ�v�2cS	!�y�]��Q�&�VL`��U�F�HĨ{�e,Ʒ �aB�m�ұw�un��c�_./��.����2/vĹyK_; _�{'��'��s$0�0��-i�o�: ����&hvU�D~�@~q�\o_��ӓ3�u X���ҒPU�$k���ۮܼ������5�}.��`z�Y'mTJ�-"��[ '��:��+�����|9ߗ�l߱ٴ��JJ��T��x�2k�J, bs��W��1�8Q,.£�0��RR�`��hl#l��1 ya��=W'��Ջ�A��H�쭂-�G�|}�;�@](ɐ�9�	�Dz�iB5��&뻪"�cWӨ/-�>#	� ��E���@>y���o� SO�e��2���D`��|A�c�6 7buRp"�����DǦ�@ں{{�&��q<��ѣ�~����[ׯ_�B^Z�-�b	&x����O�m�4!���CD�`" �-.��F5�a�B��j-O$㰢�F܆[����U�U�<-���8?6t��A�SsB<�L Ħ�!�P�'��Qf��-���R�tl@$�d])��ݗ_�d6Fks����]��D,(Z@)e�V�b	���N��_6/0a�xg�����.aEc�>K��D'�Lf�����ЦIJ+TgV�4E3 ]��{��+�������a$����Α�I�#���i�UT�rLC�F�����װT�!����+:n��I�Җ�V�����&��*���$8�:�I(�D��l�mו�kА�9�2�o?���ga�#��hۯz~xtlbb�_;G����k׮o��;���� 4��ٙ���kvv�rl�C4)3J�R.��&�d�A�Ț�U��D598����˽���1	� U����\�����
1����,]�^9�Ƶ'�]�1VD�.�E�p��^��t<+8��t������S@���
;Q ���j �=]7゘�fah�Y�������Q��zzz����ٙ�����[��=}�,2��G �ir�	����6��k�_�d �����E~lz�Z��I����`�N�<u�ر�-W�W������t����D"<�Lc�����,�pp���NU�� �� yg<��j�� �c�Ԁb1<�,R�uj���R�
�u��A�BUV�{za�^�:��ԩS�"ur,���uh�Ji�"�.�Sw�QT5���V����r,,[�P�gBME�v�����f,.O�E�@����\�ݎ�G�~q�P;#��|���G���-ɑ�k��X���b.��2�eVa�z�{awV�.~���};�^=0=>Ot0l���xv��jI*N.�p��a�J�,�*�*%���[��6_,YFU��D|���j��Ǹ���~�w~M�G}�MG���i-ܕ"��~�s�� h'ԫ�T<�n���cǻ{_J�6��x���z��cA�^ZM���[��=~��G��u�db0�-�P�	��[˼��*�BI��x�Z�ͭ^�N����|6���T+߰\����3}y��?��n۲��ʅ�ӛ6�s�	A���.��8��r�Pcc�>y�j_�b�>�+���K 4 ٧4�89'+*����a�Z�ཷ��w\8���Ȉ��T/���s9�����
��2���c%��-�;3��u6�۰n��-����$�4����][��rݺu�<{��ű�B�*k��D�ǰ����[�����,��R�����ɒ�k��L.�uS���S�e��`�cف�n)^uõ��كO?z!�|�F}���Y覵\�R�-� %���TQH]r�.-��������<��/6k�ex��D6�V9�]�n���ܿv��=�X�T����	���|��}<`����ARDK8��d����hAp+^��l?:��&l����U���2Lt���X���s����=��#Źy�H���h��Y��""�ǎY�#�
/J�>
�M�TF����< �!o�j֓�����,L� ���d"Օ��ƒ]]]��ds�x"UkX��~��/��W?��#j���,R!����7�H ��>��2��0��e��D`Y��*�$�B�A�C�	B�z����z�@]�Qd��`�"PI�a=,@Y�޲Fcnl��Xp��|B������"'	RE>&6�	z6g��u	��f3�|�(�2v#�Om�bs��۟���1�>i�>�w`޴��s�ڼ�p!�� `\�0���M61���SJI/���"jk%d��z9Q�ES<�ۺ��?���6L].���	�`��E��3�����0]���=��c�,-���� �csp�DDD�V!�dJPK ��ts�C����,&Db�> i�<@FpX@�x�$�zq��h���͚��CAKt\��[׬�85��W���?4"�b0G�Y�y��B�t�#<Ӎ[��]���o=r��/�0::�lb>6<���\�������0`Vx?�I�O���Vm�;==��K�����cK���ڞ��P��A{.\�oE��=�-�!+��ۧ�
�
Tڮ�g��"���y"o[��R��a�Iq�2�$�ۨ��z�DO1����Q��{��0~����曀? M���z�<����/��?,..�X�Fv"����ql{��ˉ�yɒтPL�A�s�֠&b���#x��k���X�~۶�WIS)/�g1�I������p�\8a�Z���]=�p�T� ~�T*��ᖉx)�5Јo��b��m�,�w�t6�L����P>|&m� ���k�&	&ȥ���n޶�ꫯ޹m;�ƹ��3g�����y��ө$v8m�D�E��T������끝N��0�S���|qlx����VS�i���4ɒ�*j	-�����%��[{O*"���M0ޣ"���q����,:�dY.tv�N����ח���ڵ�iU�ܺ^�5p�ݼq��k����N�>s���y!�':yn�t�cI�kHsWڅw0_K�9!`I�Q��H�[a�)���;�z}h��b��1-��
uU�5�KIʧ?������~t�S���Ӯ����+bj��_75.� �
,�� �r�����U��� 	=��][�]�g������|�Z���\�f�u��P�N>�菚&�Ju:F���m9�i�o���0�U
��su�ɥS��^E���f:���zeɴ���v����[>�[ϝ��"+��LX.2��E<G�Gd�@G=ջ����d%���oK���CNX�M���-�eǱ�v�e�;��s���Z��_�z��^ӭH��+<����<�2o��}�!5#p"�L���V02:��K���6�d�9U?.Iq&^�K==����F��{�P��׬Y�6q�˭`�@O��f#@�<O�%�%fz�X����b�ܸq����s�̋aL��RV��%�:����R#_��KҠ�V�&D*�˹��r�
CʪQ*�l3�x����j����O��s���?}����Q5��RZGg� Ƀ6oްutd���i�:�!
�	 �dQ�D�5�SE��(��/�e=Ӑyk���q!V�c-,���E2�&�k����t6�a��Bg.qzlbDC�
\�"F:�W���ϫ4�ȇ����z�T.�%c#qIN؜���&�^���a�*m[�i��*s>l��L�y9�]?�uaa!��&�R�6 �b���D�-�	�B�+�8�R(E���u��;mu�2J�1Iӹ�TL�^ +@<��\x�&�-�VF�q�@�u�&<Y%�mEZ`�j\GOW�����X!�Kv���Cd�s9�ʄqK�l���D�� -�ȸ�Q�L�r��DQP3q9�`㊘V=Y%��`� IH`Jj���%.tP�;�I�Kx�d�y�t�z�qZ�12ICNDXM�1��d.�@�����f_B���t��ːK��0�j���ec�&w,��#/������XL�y͇Ic���iq�r�jY�$��*�J��ŅT"Β�M�:dU�a�YO��m�D��n1KK،�3�p����d�u&��ϗ>˻������� J$%jDR3*B�ܘU��/��n��b�?0��*B���I��@����ޔw���<���{����� E�(bX� ��d�w߽�|�1�QU9�7a�:V$I��X�wUY�UKHo|�;�2�T1_Q���2d �ju� �D�(�f:5:6�B��H�SO=����_����3� �S#�BQ��8055s��7n *-ol����۷�T*�����+���7aͧ��>�䓅B,(�L���#�=�٨]�z~U��>�ʱ�����S����햌��EQ���]��{�o/����+4��@���ݫ)����T:W�7�W�^�+�|�࿹c������$l�������	���_|�'���H�if`���w^~���=џH�"x����kE!DB�Q �V�ʨ�$�����D���ᓏ2��2	L"�
 4�-��O�_\D}����� ��À���r��#�}���
��1Z G��h3��z�kkk���s��+T����Ak� ��z�>s>Y�=v���~�#��{�?22��7�C��:�.�tbI��:�<S;�04��D��R;2��r�T���Z�W�]�l�sD��s�4�x:�!)v&}�`پ�L�����J��ᗱ{~���dA�K�n}��Z��)]W._�xl8���UK�bΜࠨ�C;O<v��^�����\]-NO�>/�)��}X�t��`y���"#ɂ�/-��kq1_x�Y}8s�����F���q;��|�t����}���o���/�}6o�ٜ5	� x��(Z�O?�}�Ж��J�H��}'�qcՍ���|�������li�顑�X��n6�O�i����}�̅+��$ǧ�U�,�{���}��}?p\}a�
�X��vz�˒Q��a�G�Kk�yQ1ǧ&v�<�����k����ueee��=������#��$�ò[�E��ģ��z H��q����$�N�Xo��VJ�f�4�}���I�/��˷n-�����UN5��,�1Z�E<���>��A�m8/$��P��9�Sn�/3°�g�2١���Z>uY���~����Wև�Gc�����d�$ߏ��Ѣ4�x�:(&`QՀ\�,�t���n�/���P�4��(i�'lV�`-��_�1719���Z3��'��oq�$&Ө/�oM:�b�BAω	E7޿t���w��#O��]{W�V�0��/�O��+�������� Y��>�4�r�0�M%����ҮܐF�%����@=��%��`�������c�L¼�v*ѫ�:���0b�l��Ϧ�N/_8�q��見|�eE�1�&�3���|8��D�!�,/)F���JÊX��Npp5~����j,,޺z��!q3�NNN񢜄p��ѱ) Ɔi�	}�l�G�Yh��}�a8f�Eі��0ٮC���FÔ X�L3�:`��J�*�X���Py��rX���ӽ|��o[?*��f��z�,���
�`�V�nݸ6�Q��C�$��������u{�5�v����#�h�v��p�J1͙���h��+�v�ee4�����Dg ����L�A�]���Yx6pC^�<I��,,h�,6,mPfT|�k+�`:E�0����t�OG(�!-72�Wޱ{@ZPr�� <���ۿ��ϱ	����������"�O>���f�H��|$ݸrL������ܷ���x��3åbJ���O��kd������F>��f�p%��v������w�ݽo��#�Ç}�00����ad�@�32\*�< ��d9������Ux.;w��	�ihX%��O<Z)i(� ��߱s2�1,��˫��A����ɓ ��]�������`�0��TU��}���F���.!��詩����r��y�GF�'�)��
(��ݧ�~n�����/^�HsAt�*�ۛs�U;��g{�m8�	�A���t�]D��Dw�b��ێ+w����.,�/~�?�9�|pnCc�N�R��vjm����+W�|�����k8\�Z8��^�tΞ=[htb���Ȋ���]�?�!l�CS�1*�R���{OH�~3�m�Q��YƲ=�yZK���+Ȝg��ַ_z�;f&��I���`���ޫ��n�c�Fnbrl��L6�w<� GG��c�gߡ]�����W��RPUq0#�4���.^��Y�҇�ܮ�N���{RZ�L��k[/��{��s��}��_�җ����O������q��:`Lh]͎��PS���5(o�w�-0;�����v7J�L�|��'��W�����Iߑ�f�0�O�c���1�Q����o���/b~Ūqt-s���n	ɇ�RI��<o�7���e0�
�_U̘���PR�k�o�G��v̱K����k�z.���R9�=�uI���|����I�X��U�ѪG�'0,�� �z��F}��'"���rx��Ud؀Kܘ��/�^������'wN_��m��ӣ��gsC�#?���nݸ� ��vB&V����ݍ%���~��ق�,�U�pi�W�#%÷<~uE��5�c�[Μ�_\����X��������x��եDz�S�:��%�c;K_,����wn���,���a��,��\[J�9�k���]�;�b1;�E��7޼��;�FX�ǫ)V卼�W͊��H,N9%DǕ���5,bC�ڗ�i�B����P�ҭ���J`�mV��a�և�gF��痗��[?����r�'�z1z~,����=�.N{{�O��0C-ET2�|(��˫���h:�_n�dn#�.��W�X�X[���4G�D	_�yÈ}&L|Y�C�����%&@9�mu��Ri�z��*��vUY7{��(�N]�ע$�5��X�ݩt,-Sdx�V�NO��G0`f�h��De&�:�d�D"��5� �L�( E�z�vO���_�_=f��~�3�1�����f{m��2�Fs�������vث��np�x۳݆�a9R�'D�dk���U�I[D$�λ[����r���������n|r|�l�Ja���0찊#�����:Ɓ��v��  ץ�9���1��(Ǘ9vfv߱G����|�������CƧI�h�L��g� ��!�d���|J����a��"L�\���$�	4E�qu����T!S4ә/i���X��"OÆ8�*�`P,�EQL��=H{3 �Џ4C�P��;)�IMVsY=m�1zEԘЂ��b����#�r�à�:�����ի�dln��]�Ҋ�5�'�a�����L�k[�t1��GX%�x��6�b�滗�6��#Q��f���Llv6�P&�]ݘ�%����û�3����M{>�Kzҫ��&@��t6���qv�rC�dH'Ћ��P �5Q �H�����a� �ڪe�P���>�X��%B�)��e�6��g��8�H��a��e��$���3y5N\x����-^�x��7$��Y!��X�.�V���fTD�i]��˗�"+K�O��nv��q���8J�2�nޮ�+��=����+NX束����Ȱ2"Ξ�5Mr�N�Ć�yβ��|lÁ6t,��f:�)VVW�V���ɿ����?I:J
�h$I�7*
�h�
��U��>�~\G��Ƅ(��R�V��Ҵ>��|6�n6�Z�e?^��"i���!]̛�ܭ����S�߿zz@g.[d����W ��=a�P�'N�ݻ���ӨD�ʎp�#�m�8�o��0�$8�s�#f�Po�M��x:�mۜ�8I���A�)���#eb��C}������u�%�|���}"�t�5�211"�i�,��drZ>W�xy��N�<9�cjvvO�L�I�2�v{bb�H��e᧴F�{���<	��H+UU����,h���N#�yp׽���P�g�0�D20��BMdF��}/������l��G�p���W�\�t�,�iS*hEFE˛͟����z���O}�S#c#��:3��T,�th�Ϧ^ᡠn;�z�_+7���oޚo4̖������� \s+&�g��|�4�f_�~�?����������Eؙ��:�E:���uOH�-G$U�,8۽���/v[6���萦�+���rec���1��,t�^�T7��6� �f� i4��Q۬�j	��u���O����sJu���D�^e��|��3B?U1N]*����!xu����᮳�+XN�i�`;.�X�~�u��uΐr鬢)q���
���]�؃��A$��b�^��g|N�@�5,[Ỉ��{�9EZ�t���(kp�o^��i�����ia�(�٨`"�C1��QM��QF �)��>y2= �4��ы�T��xs��R_�mQ�IH_�u�V�T+uU-�Z*�LY�+�K�Zi���Bn������ .Xk�3f���c~,�;50PQ�}�V/��v��9v�Y��Cþ���c7�Б"��9�,�/���K�X����A��p��$0�h��|����A��`&\�I��y��{�j���#�T(J Q"^5��	�v� Jg�����w��y�t«��j �f�u��-լcl< )@ֿbSJ�u�N�PiX�Ӟ�̟6R��2Xy5�i�P��0����2x���4�Q�j =�-?�l�S�&5��յ2`�L� \ay 񚢠:�RC�;Hd������B�H��-��-���}Ya45y���7犅�L��;5���l�[^]���GB�� ��=��#J�|@uQ��E���Bb�2�1Q�y.���s�~��� y���*���-��)S�=��B� �%ճ-����������4Ul@�$Q�aO��~��ß��?~��ko��F ��	n#����{qq���ex���O�� l�� @�%�f��=k}Tb��TDAq��ʕ��}MQS�=����=33����'
^� �	�l��
�$��}�3�Jn�(��0�P1l=If
��i���v��JG,*9�p�a�}E�$JdM��F{�ʥv
�ahl\ͤq�b�ȊB�؍�J�ՕM�*18s&�+��������
���=�$C��؋�}2,��&g�Ƀ�SÅD`}NRƆ�b�/�`h�z���,��>�`�`�$�2� ��%�о���zl9`�333c�1��(2��N�P����͵�(��k��4�W��Ji��ooϸ�'}8D>U�״���<X��dM�_(���S�m`��"H��F�^��u�O=�������6J����貚����r��L2m��V�򜶡�����2�'A�`a�dc�&%2�"E"'�^��ңȳ{�����'��?�������}4ݬV�Du��f�Y�_����_����m@W@����677%I̐��ѭuHEߵ����AzCp%��"���G}(ʫ��
o7�nc8��s}�>��5�h@ ��������ܱcGG`p]�ơC2Je�1�5G�3���4�ʶ]�d��]Z�{�����?�!�Ai v�ܝ��wڠHy�D#KD&�ms�I�ܵ����h*V��^�\C��BJx�V��Bd@t��]׿r�J�՜����p�b:��d�2l�b��@�px�"��QD҈ols��Qggg�Y�
�3
e���w~�r���qH&�R)����?}�Ǫ��o~�7�|;c�<v���}i�<�j�6�+��4��w�}��7~<<җKA�p��k^^Y;}����T&�m�M r <Z��s�(�F�f�h��B��B@',ˢ���������1���s\0�T�����G�^���/�������G�?�����mc�X�RT�>w���0���1g�!Xs8�p�����|:f�V�)+��O?Ym@D��5�_��}�G�Ǻ����z�����3��(&*;�"�Ѩ�9����������Ǡ�?ٲj���O�՛]CϦ5�v`wF�2��w����r���[�6�'*����5JCQ���!lL'`1�=!)(�`Ҟ~��{��v�"��+�L]�Ñ���v�M�(qܔ����]�E�������f��"ۺ=2��k�ɰ�Am���9�`\c�{a�q.L�uAR{]�Vs=��gۗt5�\�n	j�2�$�
���q4��lW�&��0�����n����(؋39�̔Ĝ�'^�f����!��,*s�u�62"�H.���w#G���A?'s?A����b/@-2Yʘ�%�H��sb	���K��fqrOdy>�)Ec
CiQF�/J|ң��"!�~鏷XFAw�Scϵ3�Ι\���61��8t��hM�"��Ve"(�&0���bIf��ܯ� (^�&N�nw��)��`�U�5��o�6�tC����E��Y/`B? Z��>I���*�Ew�ŭT*l�f�Q���{���������J�tC��ʙ�;�	��ma���΅�vK�%%@�����e�###�ry{�a��t�d�6��-�5]��6*�8�x�����خ�����������5�<iEN�r"7�s�?���虹�տ�˿����Y��-�8U�v|/�c��U��0�c(��0eI[Y���}��-Y������a�-��23�?�ч:�. ���͍�{��k;��� ���
��ܤ���B�-9��M�Ŭ����K���a����@�L ��3p��9@1=��ܳ#���58|�ɱ��V3c���	���kd�F.���V1"-kN��լt����OMr��Eqȱj6S�1��Ꙝ�����Rvi�_���w��a� �V%d;A�3a��;iM����@Q��ﺊ��)e�`�[�cs3 �ѡa�|�,\��(.�͚ۋ����}�w���(Wr�eh�8��*@�Ҵ'C�~�>����b�Mb��gF�fg���볡��z�F1m?��ȳ�LM�x��˛�����j�����}��˫�:C&���eb+�6/��ƒ����3�4=���hU�ʹ��knT�e!Jkܟ����#'�L����Hn�:Qil����Q�������hp��CxN�1)g�_��~\1"bwQI��PW�^x�����/g2�O|���Ǐ뺁�QQHY�(��R%�F����T���y�N�� ��13-�2�v��uxY���(�J`�1Q��m	�K��Q��l/u�K�`{��*�����'��"� �:�ܫ�qכޙ��?���Dpw`�dU��1.*��
�)3_*:|��Yn6k�.�S��D��%���:�o*��%Jp�o��tH�k���1���ɇ���tr]M��M�7`����~����8=6s�ȱ�zX�c2�9<\_@�~�L�ę�X��u�hre�Z��Ł�A�
~��B��c��"���+��d�,�ʅ��R��0&��ۃ 9��#�+������(���c��w�y+eh���H D�	�� k*��u�"�y��c傤J�W�>7{�l:�<��	³O?��G�����ufM����奥����g�y.[qz�L�c��_���D����p�h��>���Lѯ��^�{�� �דYWR(��X,��&�ؗ'��3I(I1��d�_���$�� ��p6� �t[S��f�0�.� �.�ؔ��<�ͪ�wb�n�^[]�V� ҁ
�m�j誜��*ZӮ;v; �z�'0G"� ��j���dk@'��%"�i�I��@�&�&�����q�v��S��pm�0�y��]�� <�n9���d�V��A4w�4)S�;�a��L��SJhG��D�)Q���V�r�V�Zˋ6����822\Y�P
�Z��# q���5�hqK:yDJ8익]��j����\���q{n�]g����.�i`��es���,>����+��PyA�0(���P��rc%p9ߍ/�C~�
���x8������LF%��a51=ˣ]��PnKɚ'��>�&�.�k�j%(˻w����_�|Ϊv��:�Q�'�02 [��
���E8u�}�|�����-�
y�""�9�j���a���f5�ン�s١�s�+�(����횜Rggg��Je	X��cP�<�.�*�x<헜G���,=�g�G�s�$b�x"�R���c�/��=ng� ]�C�M&�V1�4���M�i��� Z^Y�7��$��9�����x9^�v��o���z��ެ�n\�����'c��p�Ţ�8(�X��2f�٬�����jZ�����B��9u��X5 ��=vb����)��w�8�7���/�뱉�z�}�܅��u*~�=
G3�Qr���pˢ$Y���X����^�@�9�M�3k�d���E��h�ւL�B��Y���94қ��/���.
#L�p\vd$���F�&a�R˨v�:�뽮�����(X'�)U�f��!)��8����tY����T�b1!�!�!���1|�������}	,����?��"�T�I'�e@�Y*�e�M~�� ����g9e�U������-�0!)^�Ca�� ���(�euv�d���v�?�Gn�Z�-1��s���~r��ś+�D>�P	�S/~������S�eryET�i�:V��y��3�B˲E.���������omlTY�zn�^�5��`*?�B�9F�=�a%mt&׶ݣG���\]Q�777i&��I@�6�뾊�?����~ރ#�4�N�ww������ɓ'����z��K������qg���CCC��q6���OE��۪O�7�����B�橬�]�L�]�w�8�vŅAa{!�]J���-��Q�m� �d)M�� ?��KK�� �^q!�x,,���d��ZXX�yv����q*�M/ɲ�7n,,,�
�b�`�qX�,OLL����r��x@�q��}�AS��Y���8��m�#/ٽkǞ]{�V�C!�YN�ۀ�k4��fhcvv���ezG�����d�&]@:�v��9`*(]�cUi�][Xɵ�5 BTJL	uǔ���;��J�����'���E��<0�j���믧��#G`�y��CDӪ��t@���MN6��D��/Ɛ��l��^���eQعs��i��J,�?<��v�?j��M5���Z�l�>w�v�4�u�̿"D7�]���F���}@ �vJ�����yZ���*��L:��պ�僅���4�B�Edc�ĭ^[5��fM�ġ��mL9J�E��)���L������r�$����B��ھ��0r���X9��E��Y[Z�Z��kN���f^Q=�!H����]�U4��S��H��Dd�*��١�&ݶ�ؒ���MUJ�Z��\[.oF���\�Rl������;�h<���EOX�JW{��&+z:���{jb)"o�ȳ�����j;�HɖB>���B�%| vW����E�z	-}"oH[\�D�* "�?��{�  !��vU���*�,�x��4���r��0��Z!�c�
��Zm��lԳ��!I>,�AE��hK� �ȏ��޸z��VR�V�M���	�a7+��D��U2�
� �ĵl���;J=-K��\@X<�gӀ-���N��լY�qxX�ƻ�U�lٵ� �([Ra��깛U�Hf"�'����Cb���)KQ�eຂ�W�"?˶;�n�ڨ-^K�����\�Y�5�k�����<g�jt�
��%1ųF^wY�T�3ɽժ4��"Dˉ�̾-
���\߃�Q|�����q�(��S0��GUH	������jݺ5�hݜ�
P����I˲�W�]:}��?�v��]z�xz��+W�� ��\��UF��;�S%����a;=����t���Q��}{ʕ�f��i��4��lnR�x�ȼ��W_�ޅv��lwZ?���p��;|!�ڗ�f�4Yr?�	�e��x��zce}cdf
[��@Qee�T(Ć��IX�]B:� �DK��sZ1Kjf�H�IVa��\��X���	!/��U�[�r��l�@[ � r�P)��ȧ�SP� D�mY��$H�<�P��K��!>X%�±a<�=���)"/�5�~&r���eHRz*?>Y*�8���?(�P$U�음���C���_����Pa������1�5)�#�T�ɹ
���h�'��`dsj�q�����Jn}�䎕�-{cU�:`f��կ��ɤs�����v<KU�(��Y��}Y H#����ޥ���U_-G!ᇔ$N�M��B�ĄZ�^��`�Ǻh/Ǫ8��W"�bs"!� (��n�w�L!�3\�܈%:e�W`�?���S&]�� G:��*(+L�Y2�٦`e3Xr�C^�t$Ӽ��F�Zv��i��,�s� �o:L����:C��.E��g�2w��N~h\��a��6�n�� ��^���?�����Y#�*āmk���N7!R҉���T���]KӍ���t.�&�t`����tt),N>��J��NV�gY����#p�*�Tn+K���#��C�=v�V����:^���>x萛���&j�j�Z�cc�ڭ.](�g*�rm��TJW��v����ZXz�&
C���#����x (�}�O�v項ڞ��
���B�Q�;�Fyc�u���������5`�'N����;�$�Q��P�#p�������2-�֙L���v�~���ru}jf�dHU9ۑ������`���9A�!�q�I�/'�"0w����<�߱��/��[���N|��Q��ӳ<a�kU��Scc�>u"��y����^������rm�n,/r!%�c�Cn2���w�q�@h�Ū�(��������;-��kimѷ܌j�;�kbׄn�=���������/ܺ�|#��,ɲ �dhd_q_9����R���!ʀ2Qp�$E%`]Q`�z����|ab��gǡ�q �0a�n4�y���wac�bvI�.�	O��Y��(5�i[��F8�$�E>�+r6b��o�)�15�wdJR����Tٍ�f��rku�^ިl�  ���fAd�. E��^϶�0 ���WR�M2B���
u�X ��p�[Տ��5>3��4�X������7�.�?7���f�%�ݦ��n��^�����=��{တ�g��"`9@�cYJV.Ǣ��莃+):v����y�z��ť��f�fT�q��g��P�`�
������4��tܰ�n-W+1ό��||����]��b9���ʵss�s��^u]3Gdl[�>�%!�'��E�<a�[�F���AL3� ==��n������w�֭[�Nsx8����ѡ��X���嬯W6�+^�"1EI�p�u:Ɓ����ТQd#���'���� 1i� (�Ĳ(4�83q+��F$m`���H^�_#7�	���(X�D���Y3��xH�^���� ���Ï5[����6Qׂ��,�\z�e� �����L:�o��v�����6�t*'�(���O_�����촁 �g��)gT6�6y.H�d���g.�=wCUR�Ex�k�K����\�
dǻ��2t���U�J�%2M�Cz�|?����J�k��4��Qp���!NA�r��������X��2�+q�,6���60Ϙ��-9K���,��1"�q��U0�j��>��KQ"��;�d�tCҵ@�D::��4b������`]��PR%�ʯh�܎X��v&�0Z`C��!�)L^�0x�-�ab1c�dY����O���͖���)� �C�&I�@r�a�vP��h�`�z�d;���A|��߇'i.��h�a�J�����8�%bS<|��ȎY/���S48�����_��*
�F}<��~���'Uv�`uu����^��fN%@�����v� *�|��bC@BQ�����y��O~�CS��G��n���;{��ѣGC%�Þj��ö����_\>r�2]G�>��׮]��!���z���A~`Ӽ�kt,�c�mm�+�W529~������r��b
6���Đ�����e0#��({�*��%'T6k�����Z�4�"�K��hԟ4�D�c��}��:�V��!���?���M��OV���íI�b@���M��Zш"�AF��>��6�b�Iz���m�%L���������ٚ�����QY[�i�{.R�(���Noym5[�"7�Y:�~CA�����������cm�����kk�P�����+���h�6���cd@v�ZGqD���^��+��<1>:� .C@ =��Y-�'�Ԧ�
�� ��IW5�H��\�C��pl8��f�N��vH�ON���?Mьq�׭7����r@��9L��	=$�<��4D�E� 
)��Mn��/��.\��c�|!�V-�1�78�X��9�Mc)Ǩ��1Y����1�1ӓS�tb�٨T�˵��UC5�%�ǂO�$)Wkk�J��$Q)����~�D���)Z�!B�J��#��%�|W�Sm6xUN���+W�^����'�س�N�R��a�D�rۣ�ӻ��g[��F��t;�BEc����7����I$��P�B�I��ӵ=ߎ�|�85��116�gOqfZHz�8O} ��X�>��k�{����טHd�G.��0���R:ϐH�O:y�X�_9����Y����w>��sǎ>82�cd5L8A"�	�fd�ba(��k��6����s�nXwb
��>	H����B���P�6�p�0�+(pܥ�ժ�?z��O|���n���&�8�%
�����[��y�'W�7�v�˪�j��K
B��p?&Ql�e6ĶT�=�Ly�0����A[F��`۽��=rd�^�0ɨi��b�9��w�����+?~���J����r)�E��$ʰx!�M�jl����$!˅���F]��G;����&g�H�,������{���Б[O����/����M��ђ��I�Kz#p��}� \`Ŕ�U,wi~�8Yz�ǟx����]��	����n���ד��o,��ڀ��TIOhY�ΰ.~��Ʉ6D�Q���P*�V ���k���"��up���x� ����� ��ū�o]�ڨ9�N�E�6p�� 갼+H��H��xp��x�*�2���24����`y!������/9Lt�nB{��ڱ(���C�eE����^ؚɍ�P�c����9{��o|���T�U�4#| ymc}lr4ef�?��s�
#�NXZn��p���۝��z�w]MQꢂ�&Aw��<�Ѕ��h1m�"'������"=�x�\^#P<Pd!��0�s0)G��WU��Pt�c�S*��|lC�:�q�`s�|k��잝@�,�6err���z}��L��֔���XU���&D�#
I'8���_ B�1|�u_�4.F2/����cc|��(�x���@�	e�\J<U,&l�'L�)���N1'�����e�/C=��8�ڋ%� "�HTٰ�q<������xb���6��\Z����r0)EY޶in��,p4-�J�6��.�B�{ݯS��z�D�Pa!p>/�9�=�)'O��,*'��;fg9s8�8C6T�� q��Q����T��3�߱w���aV��W����g�F��)�lUWC"#���]��`)VVV������={ga��!bϝ����ҷ�~�֥�G|�������t����W��|�<��"�s��~���� 	A�Ǹ/MZ���j�w�%��`�_D1������/7��?��?{��� ��U�|��5 ����=s��ŋ��ñ*�
9�vOmss�^�W*���U�s��<����0��,`�.��݄�__�~��I#�q��-��ȭa�	�Sb�W&<7"D����$UB�E8�n��۸F84����`���l�*��*��	Ime�x�u;@�B�/D6g��v:���k�v����\	p߾=ã��6��4Z�ӧ�V����;w��RY���0(� I*`r\ ���c}}}aaicc�v�	"��S�XR��	�}���l?������3ˋK�ӻ�v�赱�	�Oe~x��kz6�΂a��V!kf�Q�@i꛺�2�g�8C�*9�il,Ї~{sLz��nu��IB?����#��
T��W���	�t
l̊	��2�i������˛�����ʏ~��SO<L0	��y��/p�E�B�����K<N�a�;˱����dJ�R"!���>�(�w����4-c�|�Z������B�I�q���)���2��02fϳ�77���,��?�����灝7��O�@,� �$&Q��mL{�Y û�]�'G�y����%[�T��P5X���	0���^]XY��ҡ��8qt�X$�aL�)�s`�8-�y<ЙnT��{�0~.�p %x�c"Nt�~i5���B>�`��J ��V�R�����G�>i���(t�����6�/�����a�T{_��wz�*�O(Z
�U.f�P����k��m�h	��$s���Ԫ7n�/?������/>p� ~xq��Jb(j��|zh���P����s��v#M`$��F�Ъ<r�я��9����Sń�� � �`q�;��g����wL�����D���L��N�l���
8��;��k;�Rd�X5�f��(�s�-�/7ǂ**��ca^���Օ����}��Ώ��\�b6r��"
B��)�3Ie7�X�N�Z��C`$��%�∦�^���q=[#��l�u�x��O���㓡�݌�\�j���Ƶق�o���˿�ʥ�5QʐV��<�m�D_��h��" �~I ��hny�ܼ17���>��?���rcìl��0t�Xӱ$ΰv=���o�q�ӗ����n���MA�T��\&�*3�Tw�?*��q�'�T�a����1�鑂��%�Y��D��d�M� �OI��$��Qg��N�{���~��[��H�٩��ƺTk �nwj���Z^��kv�&5��ewQ��q�-�w��U��8Zڿ��$�
�6ؖ�;l`�+x� `s*�b��k�޶����fk�#�
¤I%>X�4pɖ� ��,�X����Z03��LǱ��]o^��X];��gƉQB�H�`l��w�OВD!6c�DT��YW��^�T�����,���ǰ�ˊi!�QE�$��`N�#�H�0�5��P�(��Ӑ�tV^�#�KT�v H�|?�=2o�����c�0�I��[�(�� �_�{�v��L+8nm+T:f����46<44�[���A�Ǡ~i��}lu�c�,*����܁I����Y��"���v�=(�<#+	��}��� �cš������^��Z���"![b15/��
�<ϧSC:��=GĶ��Gy��^ �@lr/ʛ^�v�?�O��rWS;��W�7n��v�]�p�,0�#GOf�y0㍞U�����O�".�3)]7�毓�Q"Dhsq�p���=�UT�$�������k?:}�̱��aq�ZI�e	;�`��@�f{nn�ҥK�N�ZYY#]v82�V4�P=�#��[�=��(�������Ͽ��;+++���Z��d	�~��wk��O9\ޠ�gP7x��Y�L�L�ʩo���밋�`��vi�c�]��j40A~�%tt�h���~��ᵫK׮/�������G�>���|�X^[�z�,ߥ˗�~������aڣ���x�����m#)�3M�
=���?��n_8�{�����'��w��[X!Ib�
Em�Q�i^,<c9��zVw����D%��A�N�>V�ƍ�FM���	����ln�%�0��e�TU���7*�F�V�u����]��
2Do�Z�G7 M�_��J�<�LҢؾ �JExMU�H� �驥��յx�bN�u�r���F�(@�>������P�cY^Y]�׫��U�5�j����Ș�g��
ܣ�پ�K�մ6�+�U������. c�/���#��h0��Nq��R̝�j���h�ez~��ҹ�� ~�}��2c�7Q�n��Q��^�U��D.Χt�^��w�����O� Ќf7E%�2&�W�WnF~k<o>�я����u&  �h%l�0vc*[$b��� :����w�f�g%���q�f�����'�zad��[�Z'��T,%mk�Ţ|��d��'�Od���W��L�^M��&���q�Їm�( �Xdc�	ςg�0N\��w�F�T���O���x��q${.��!�`��� /qk��*����>��*_{��յ��S\��15M�1�u��.`%0�[Ek$YL�n ��zvhh��^(�������k��=?pb]VClX��
Fa�ȃϹL��S���c9>�Ɇ�;A�
�7��PY���b�� ��H��eCc�\���t8ᣟ���́v��6�Ṋ ��1�ծ��k�c�{
��3��o�Vm���[�2�յL]� 9�qP�P8��.����}�o�0���펤d4^S��k�x��y�ȍ��Z���m���f��ɉ"y�ב^{�1�-�>����\��I�x!�}�P��j���d'{�8z��9a��㳟��g��"��e#�<���j�O�1F&N>��V�������cl��Z�ز�(�!<>�� %
}Z{�!j��Is��Bb����Pf4�TVo<|�������L��m,�i3��� �V-�A�d��ك�s��w���C��퇱�� ����/i����=�Q*�b��2�y!��$]a�e��3�^�vm.3	�~]�׆s�0�%��X�Ϲ���'l�Ri!��A�	_�D�n�s�㛇d�+U1	��j��?f
���2+�q�V���OD��m\]KEY_-ţQ�_�B9�XT�D`�Q�� ]�r
��mcQ�!�m��g$�w�3o�������l��p, 4U�Kfb���$V/��l��L����Z��Y�r*����m�6d��C��]�[��ąVYĤ�N.�cP�D�T2�5OJ}�NX@��(Q�DJ�o�6d���a�#=��9	�ڍ�~�x��dZ�����ʴ�8�v�"3���z~�uT��U��w<6P9!�}N�2H��q6W[���㏉.\S������S�/�>;=192^lٝ����雷p�p;�z�Նa�[�c�)���Ӝ�������]������J�9'y�w�g�$I�"O��OB;�%^�ŅUl�Ώ����������(Z_^c���Uk�;���㳩�D�fe
�����]�����
[P����F,�6�n�~Ć�Bm�.�\'�����Rs��O:v�s?����/��������c3;�X:d��� ͶBK۬Y$g(R]���JB�!c��ܒ��cR�����]�!}�*N2q�HH���dvvLz����Ͽ�����^�Z��L`b����*T���ja[L��q�[���o�����E4TUN5:���\*�5���F��D1����"�7Y��Pc����[cӑ���(���rA���n���x��@Yn+��'���X+�Y������2�9���ɚ��u�ȉڧpJ��������ǟx���կ~����� �07�J[!T:�
����f�/�������=��S=��D�J�����ϗ_~�\������z���Q�����"�,�\�궜^S3����b�od�C]3� �����!�[�P4��0Ǜ{��G'����x;�,?��X^����u���@��@�V�6�O����q�6���e d�T@7��M�<�m��^#l��H�Cg"�dl��j#�R��,W֧�G��y�SR�nv�����|�Uk���c�<qs~���3n?�V��i|���fjt�e��릖Ϧ#��tQ1#�W�Z�ӓsI��.3��F��*�P�R.HU�I��H��
����u���ϒ/����o]	����w_�{$�T�w?B��Sk�k��&5]���"�ZǤY������i� (WNɑe=�A=�*1��R�B/�9�d�������7�ݎ(	p��$���p��j��g?�ͤSy#$��s�N+�+>���c�6��6��\h-�o�<���ݤ����'?�>_����V|�������)
Hl��A�(T�Q��Eؙ [�|׎�|W%U��:N��Ipqж|�)�z��v���O>|���ƺ�MM��p�,a��K��e�"����v:��nV"��hv�l����w����I��e-WO��J"ֵ8A.��↮&�;�:th�7��)�59�b?tA�Ddcp.��*��	�M7
t0��L�vU-m�É��̳/��w���;U�����d1�+~bc#��n�q
����y�̹����?��s�Rq����İ�0��:��T*�<n���"Y���Uk�Z���ڷ���jn��8���ǖFp�\[je�3֮�lq׾�����7궚]I���m���f��2��5=�Aa`U{� 2���=X�L�O\����j	�T@)��~�RGN<r���wޘܠXP�5���]p��Ũ'Zp�9���>�����4�4RR�9<����������xQ�g��Zq��Z�_��^i�<X���Z�y����r*3
�Rn� ��(e�FW�����b�T���$E���`*������&Ù�\�x�Á�d���BQ���Ud��G�5E�<�6�������#�������XO��	��\���L����8��P�J����@3�כ��{����umka~����	3@脤ن�LO�V%����FR�����o-.5F�l"	�7lb��ĩ�[��
�H��a��1�>�Zuns�V�p8��N����7<_VK�9�P�M�U�''wlV�=��R�.�q��f*?4�%u6�EA#�@"Eķւ�N��'i	PB	j>�Uz�M��D�Ɵ�}�QE�������O���V��g���*�D-:�Ӳ
o�uS�� ��D�	|�����	��g5-�,hj�r��������+G:Ċ�C��i���a��NMM�J%@�kkkT<V�
$�8����.���Y��#Q���Q՝$�$f=�l~���$���]N΃�&zq��y�ʥ.�ޘ\4jV32V��Z�,r<maaw��V����x��1'.�s�!	�:������D1�Exk���ܹ{hd�¥��Z_�x^U��tmt� e�`���dE�E�S�����J&���5���.<�]�v��4E tuu�2��#S�}R��7$8�_�[����O6c�	5�f*&�u����)UU����v�n��"�n�]�u{[]"@oz��N�M��3(#սX���.K�3|��),�%H���g��lH�/ɴ��vE$� �8#�j�p˚jd�X���4:�ދαy��'��x�-������@4�N��4.�?]XX���o���K/����>���p:�w.&�WL�����P�Y ��M����y�Z�$d4�$u��������Aa��M�\__�{IgR��'{��g�}����/_�Y	�Ś_���$y\���
<x���t�!H,��>����!*wT��>7�[[z0�A��s�� K�"�ނ�1�����_��͆��Y!aҝ��Yc33;v��җ�TL���Kt�0���Rc-e���uC�D��I�Ņ��������_OF����?X5:т��00��[�{�������K����O}0���ߞm��uEP���<���R ��r��$���N��������<�O�7����$��`0� $Riʢm��z�ڕ]�+�J��\��Һ��e)ؒ��E�X��PY�%R� �@"�`r��0��o�NN���w���p�V-[�h�����|������2����
�	��M#Z�؁��g�&�������P��	���.�$�������f9�I1=�^�'}���O�`�\"���r,�u�i{N�ѽ�c5��G��?8٪^����|a��`�0�У�'�����IV� �E�d�!ڊ n�g�4<��y]��a���m����2������ܬ����LjC��s�i�	GG�W��tLR��w�[f K@�d4>C�k,JF�#g�� qr��8(���r��
PH��m�h�-NW�t�������0@[[
�����Ve� ��J�F�Ո�����険{�س|�V�o֬��?��(�w�jN�S(�9�t��&Z]n}���zCC��ӳ�v��DF��d�Z�V>���;l� �z����\�XVA!�sz@!=�gs�^4<H�&$ɼĤ��i-��I�-�G�F'�M�N��yf��Df�����*�"�r�$�b�䚣G������L�����t&���Nht����'�)^� �����dڟ�?~��z�m&�𘪤���'Ǵ(3�(���� �bDb[Q�B�!�IY]=8;{���˝���+�sŉt6�v��6:د[V�Օ��Ň���Ջ��־���E�" ���3;r���t��|��:�!Z�Q7��Ըm��f+��h���TI���p!
΃ �� �pX�ʂp������ߨ~�ML�p�К�"���[�������[����p*�^^^n�{��ӊ�<��k���x�1��0�V������7��;��J�Z)����/_�����<0�o�7w���/\+d�2�	X�6������u]Eh  @�`Ȋ.VlZ��<337�0��F��@T4XϾ��	h��7DMp�>���?����lq���80�]k�\_il^�ճ����4f��
����Y�!=ZD��/���=Tz�`�������U�2�������8��5>�BfbRE�|?b%]� Nr��Y���x;
y��Q���5@D�YN�2|B3���=uy�_}���/�o�>��cj2��Z=3��tlY�GFF���� ���0�S�#f2{!SRI�{;wBs�t���|P%�c*�5,�d��`�mj<������)X\p=���.����Vnv:.c�ڣ��n�PN&K$�'�L'K:�JQR-�&���@��P��1�R�/ia�E�1�Pe������/?�Dbvvveiygs>\M�����IE$���Tz�F�]��r��/�R�,�Q���/��|O�.�`	�	 �%? ��z��h� ���m�G-�"U���3�v$�w}omc�����N=F�qI!�}=1����e�-�rqr����H��+��Q�a�"B^<�10a-7��1�#2��&^���0�u"V�8�>�:H��0����J\6�n˃�� ������W��U����p�ccX�@�=fވ �Z�7��>��n�P( �>~���3g^x��	a#*�J�P�����RV�9�ۤЭ�>�������vwxz.�>/���W�ij��N���O�T�O�L����[͝Z��2`�H$����J]Ap���0K)�f��p���ڜQAz����|���Ķc�.(OSu��3�2_Q��S�u>"���rDӴ�ix5	����P~�cDIx��C)I�Z��q!jΊ2,c`Up$ucd��%P{�E��r�X#�P���ջ������C$B0;�q8qa���zGw��k׮�<yr�N�L]���{��pw����n4�������`�o0: �x˥�	��^�����
�m��L.��hq�~��Ba|&�/()ԉp��L�8I�&[�f�V)'����p�G"����,#bo����]����z:�J �;L�'�P)狍��k��j�f��Ԫ�#S��4�WY�g����R7��Tyfb���7ߨl/Y=�kJe�$.A� d��P\̎Ȏ+t�l:Y7���JZRM����N��L����ŃOtB���im�:V0UA��3z�i6v;�<#������`������Ɇ@�H�'`��O��0^h���_��̍���L�5;A$YFwk{�k��:׏�F����ёi������p�qY	TXM`��O#�}���M�H�W�۞�٩'����i��ַ}˙����2�NF��j��������3zZ�T�5Y�����|�0�L:-�^.�D� ����T�L"��z��%Ռ�Y[=M�8���[6�=�1�.\�}q~b&�/p���i	vb(h4��Fcw�U.�d�ՄG�hl�tD^��*��0`�r'�!�I�:eA��2��X�g����v�Zh�z*[Υ���V����s1�=�jU%�^�]*���a\RGO]SY��|�F�/F8E�El��I�NV�f�F8�V[�F��gl�[^�t���q��'�ВTS���I�h������*�csO>2591ש�n6�n'	୘U�P�P�(��l=�܆��C��|�p����4�����m�'B@b]4R8�O�A����^<�x��d���ıa�����t�a#ׁ�������~����rF��%1��P��)7T�O~����А�{�IŹC�?����	NU�vSQ$V��l�����t����yj��=����Oy�рu��Ӵ/0l=Ī����eq�
d.,��m��+c$�"0n۱�xҐ/��$��W*կ� e?���/0��p�Ѩ�_�ȳG�;X,1*̚�vp�=����Bj�L�5Q�Ǫ!�1ܨ��D���h#C����j�r{_T���*F��}�1�AR�5����J��	]֭V��^�0rʰX)=$�EY)���i��N�=���.�������>��G�dvu���ۨ�����ET:ݞs+̱����2�C�I�nj4&x��CB��aSv��u.衹�������?��S�Q���hwj,�3j�c���R��W�Tƨ�N�O0��a��繬��迄)���ar�����W u�����X���F�`��V/��zukk�z�� �at{����َ���X���b�U%��ƉZz,��(�ȅIOj*Z@��z:�=�/�ؔ��[If	�*Lux�3�OR_ �~�P;`1�C�˰I���������a��k�N��x�+�w!�u�@�0��vb�pV%_��
f�NjJ�"ҧF
�"�������0`b=r�}�C�w�u`��Q;�eX/�0�դi	 Ho��6�n�(W�+K��M�ѕH��7����:`k�=.\|^�L�0�8���~/Q%���1m�*�����zLv�\
l�nq�W��!/�	��I=�h�1G�N��
�m82�#N��X  ѵt���Ju�@&�胠���Q0v楓yP�<�E�=E(�E&��������А g��������˂+ H+�9�><�zu��X��`˲,�gQ�C�d:��ā�elb������ZD摆�Z��+F��ý�,~X=B���'�=�LQUa VVV^}�U�yT�1ֆ�	���|x�y����Mef��N��k��nOLs�~ý-4�N�@D��1}_�>����I7_����^x�82�S}���S|���`���*�<7�4�I��0���Oii��aCB�P�&}�-|s��y�	��(�SD�B��x���4���,����f���m-�eS�$�8F��vvj������S����R�f�����JH:���p�'��	%��%C ���C'��p�u��V�mF>g{fg����y[���lO��bη*����d�3�<�.����]MUM`xF�dRU�H��U�(�9R�V<~϶{n)�T�n\8}�����W�NON�&F�.�8m���U��C������pytmg�Ө/E_!�ɝF{(G"Q|.r��R	{�ݞ�i[���s���v3�Y�r���(Ug�L��������Q���f5a�۝�O�:qwect|"���؉Y�mO1�	�bŠkz���Ld{Fw����닰�G��lJu��l�2�j�v�][Q�`4?��5�㓚���z������#����"II����ݰ0]��Ђ�����-qWiu�D�zp_f�Z��c1��4��j�����Y?���6I"	j��꼢�Z����L�a��J�)׵�7ɱ���[���825u���K׶<FmW7ݱ,��&�Z1�(���;�k�.��+�U�uZKg���%� )����"����9�$4���y҄๙L���i�S�|	�Z�cZD�Np��͝#\�ώ��8�Ot�|ח��VC#�	��� ��|�LJ-'ԓ\&��Aʙ"�=��T:�����<v��ME)F7��*�b!1��9'd�0����W�����+�@9�e@�P L�r ד2`)�PX���@Y)ɡ.b���,�Q�ra�<߅_�z-m��]�x���@a�v�۪YV�;���PY�����s�w��#�j5�\G���"I�p��0$��M}�xf
!��H���uXU���h�!QRB/"��?)"�Lh���E�&�`2�B�9yr,%��z8�#GR4UM�9;;:�H)/�"%��R�>9=�]_�~�嗯]�Ȅ���������,���W�����+��om����'���v{<vb0�@���ш
|ł�����:�\�H1<X@>�*R�*�&d��J���a`�f�ˣ�{=�a16��e�;8Cr�����@�ıQ��z �|��j{�m�݄ʹ�d�p��47��a�s'6�O��>�`k��E<`�F���X�n���i�Y&Ĵ�n��M�2�$0������or��!��р�Y�}�z߄� �����$C�]]]���֟�5�������ޯ y���ً�{�>�0�W�V��@�vn�IǱ���,4Qߦ}�v�Ӿ���%����]ž1P���;�_�Pn�t"��I�ω#�q� ���4@F�xL�"�v=[�0������D�T*ǀ��1�Y0�q�Ս�R� �+iW| ��:%�Mq���[��]%ԓ�.@x�i�J���L���c˪B�0p����I$�RD�ّ,�*1�	�ذ��To��!zwZ]HJ�m��Q��p�܋�<�F̞�u<]�ѠCJ��ѠY|���CV0�p��)�#K�I$�4�`!��u�zG [(a��l���aK*l��bxļ� ����u2�"��R��v�711ĩZ��3�yZ������]F�7N��o���z�-�G��qF�]�o�.����wO���ڌ��\�^3E���(!��#�&
�D��4d8�8���P�5`=.5�m�;o�uf�'O}����{��ψ,����ȷ�$�Τ��j��=3<;��KW�k��zw<����-,uׅ�U�P�X�g�`�b"���3߱���o����K��}�Y��G
s��պ�(z�J�j���]����\c;����GFr�3�$����vW��&r���cB�4[rd�E���~�HI��,A�q���\qr����/���;�9|ߡd1�x2����p~�vV�\�,��c�\I�TN��:�E����B�zy(G�T��fSҳsg��Ͽ��?���Vkh�Щ5��*�G0�	1�:�����5����ӏz��?	����f�����a�;S�^��VlY��OrJ��ʫ.�zc�\z�տ��9~m��<z��g���;�(��|��U���^�|���|���Y�AǏ_}���Ry|��$I���c�F!����� �!a�Q��ó�=���W_������;p��O?��ӫEl��,φ���\�ӪU�-!`�'�u%��뀜�C%5�	B�ש2$��D�O+KCb���C�I�39q����_���o~GO-}���qqd(3�d-+�\�ezͭՋW/�^�����tVy���I-{m��nu�<�`"eˬ���#/"2	�k��9A��E�a�l���;/�ޟiue��>��%���4`2N�!�,?7=��0�W./LN��l��W|��Q)��PR�F�a��6�힇�t� ����tsrhbxx&��eܶ���ۧO��T� �%�/a��mFX�B`��a��y��}������?�	ӴO�8��;v��ٳ�N�B3��ѥ�%�N���I��^߷oߡC��\�������t��pm	�%-���3�W5���V* Ժ�V쌏c:r4mfz��݂w+泲�5v+�Z+�� ���j����B�j�z���%ҙ���(d�gg�V7.]�R.��7����n��/_;y�4�xV�E��q�����wo_\۵�����Z�9&vu���/��z�G�y��O��;\�6:Ȃ�{	���D�� �۞SA���TYZ��/#�IZ�
ga%+M�ӆ"�Q��o�i�ZV!�������^-�l�$s��ً+�����ʗ_�N�����#;�����`4�#�Z}�칋h�*��Vwu}�\�MN�Z����lَ"K�k�m��ohO.�޶_���GR��D&[Ԩ�-�K�k���9�n��[�0L>��07�/����5�������Y5��@Y�00+K2Z%<J�)��M�~Hu�Q)�$���|�C̜lۂ銚�Lt�C��c ��l
�d��Y�'�|6#����G>F`�/eT���c�F@� �e6�����+l���T}��L�*^�;��"���H�7�\�׿�� �_{��/���/\��)�q]!�=}@����nFɤN�\	q���A�w�"��'�m�˺�`:���9�eę������J"�:�0�"���������e'�>�����8�=UR�D�ك����6;t�g�H��G��ѱ�i7 ���@��
�q҃��Qh��K�|L޳��^�-�W(W� �iT��vh���̈́渨i�k��7�<����L?�Hr?VH%4�ru�&�cBo'V�υ�>�i�J��4���Ȝ���jI�g�C�QDЂ%#��g@YÀ�v"����RǱJ����Ց�U��&�=YJ���K�ga�p��L)i���A���ڵ+��5�����_w���Y�/^?@B��m��)�2�O��v'��ޖ��)S4ؑ��"� D/{D(�0����׾����jϴ6���{njl$��6��sBP#s0MU���1.��r�H�6�'�����<�G�+��fU��C>#g�k�;o�~��'�k�қ��ʋ���NS�}�D�HGٓ��Nۻ���~mt��^/B�Q#�$gxhT�j�&����pώ ���Q"�r��Q��^]��������_��ܱ���	$�g%��v��쬵�M	�^oqq�c���D��[nOT�D
m4a� �
2� ��D�#$Ax��=��%��8~��_��L1;?�|))e1rm�w�*/Dv5%�v���0�΃��Cc��^p�#v�颤K���YS��\Rg�)+d�D.c1��������Z ��I�\jvj8��`��=���U��W�\O$���o�>h�Py��=A�tE�a��_D.K���|F�9]��Ű�D++u�a���N�����d1�9���z�LI�	��ԬU�vn����,3>:�ht;ݪ�2JZ�8 C1TQ���D��a�4�Hoe���8��'��Nvf�J�B1��J�aQ�t4�Y_���oo����mv��v����)r���zz� �l�!&����}x�ٵV6�V��۴��&ܷ?��%l�`<�5N�v����LQ���=��F��OH�,��{��wO������o6�Z���F� ��!�p��Zە]��m��'4�m�9��;��}/�~X��a���
�ǳ�����|�3o��& ��/՜���v��������Bd����>��B�����ϟ?�t~~�0"8u�X�������J��V�2��s��Cש���:�v{�<<73[�W76�dQ=�5��6����aY���\.o78]���٭���?��[Y\\����[�Xmw�:����t�w���y�e��z�c(u3�%���D�yek ��n���?��gY�#%.c�3h�Ē��Ĵ6�n�$�Sݴ����'�T �G{��1P�Q���E?��g[϶�kf�m4�!:���I4>H�5��n��rͯ������l�4w7[��.c�)t#,Im����b%I���ǋ����p�h��]`A,9����E�7���\���JjPDb��/t""P��ypY)Ud�rD�
ѿ�<�|��=��Bq�^���q���X�\�46��N(1p��@
k�,����cV�z>*�5x�带��ɡ:��{h����I���N��Q6��Q�X*��J"����b�k�qSQab� _���hR%�S�ݾ!�;��,��e����u���&��Ï<���O�w._��ܞg͚�hq?�`*~��W����!����?���������Qn���w^"MD�A��M����X)��L�zF,GF�$���~����Rq��?����G/�����2�+\o��i:�J��a���20��l���v����t���d��}���~X����o��5�90�rf��S��7����r#ͮĴY�8\ݱ���IQ��:��������6�^�T��Q1����x�#!�����X&�K�s5f�!��!q�BlL |�Me'�=�v� B�]�����e��ha�>��Q�v����h�����E�� ��DU���`V�J����E5/��X�	V�h�n�Ͼˆ��C�n����\�{Ex�r���?Q?(�Qp�0�W���u����������/����h��)+p�i�@�r��r�Yo\Z�~��ڕ�����?,۫�M'1�(�"����X�����%%�s�/��o6�/��gj���n���<5]+���͕�,&3��e.+K� ��wO~w���W_0��ʇ�}����[׷7�L�������PR���ݦg�	iX^�k�t�;}��?��[ۻ�^>��O�������+��el��<`V��b���|��Ź�܁�O�/7�2^�l���3�ɔ�+�Q�m�u��Q�E��X*�o�~���lAO��L��offd,U/ee]���\��o7[Cr^_�ޮU�6�C�FGǇ�<|$U..67vv ���M�A�z�����%�gX���덍�'��7����Si�$�T�UP+4��0�iux�81;ԭ׮�������O��x���s��0����Ac�uQd�ګ��P`�Ȏ,Iӗ�v~��$��v��_����S�r��P&��I����$3�i=�r�{�cOD\�P�g����;����\�PT���9W�d�{.�E�R&r��}�k�N�:⌬?��O?��A`˞��������)�?���VN�N[ɦ9/<t߁�]����ت��\!+���G���춂��c��醾�6��+k��7�{��?��w��ᐅ#*�"�2pB RjJf9;2��e9){n;bmI���޸���yc����o��
"�qlਞL���Gl�Ӆ���̴ hp`U�0PT�[�7�0P���l����	���o��ųX鷼���r���W.�w�Vw��$:�νz��[��}N�}]�e�6�	f����W^�kڍC=��Óf��)s�.q·%�@��]��� +�smkf��acgK;4���t��P���"��	��ꏂ�>�Ax�@�@��n�I�|P�0���v�$=� ��{&���;������zY"�&�Y�rq<vL�pa$�lh�S��:ĊҎ�RP�QR�r��`��d��#�����[߮�vk�FRz [\�|]�Rdo#%2��:W�������&&�k[0- �w���F�4���aRO���N�����kf�x�F��$t�D 
�����?b��M�w"Bh�̋0�,��,�^�s7(��Z�P�n�:u����� ��c�"'��t� By�V�r�ĉ�~��i^�#��0(�~��(�����$x��r|�Re��#��2�2�"��aA����:�HWD��lon$uE�|>?z�P��f�<'~�С��m�l	{l�\���tл|��8�Jڐ�h��V�IG��,�\�O
~��3��n�+�0�o��������z:���AE�0a¸!f�{Č�&^�8+H�8|5;���bޙ9�E�I!���$�HT[I+ y�ʨ�Ija�����;�b��@|Ϩ;�^��v��FFF�Ʀ�{��7ϝ?�{V�,� �ݦ�1��-�U[�+��(h�'n���(��߂�\�_C����0~X��e�e�0-� ��U�D� I���h�O6S&C�sh�m�r:�T�-������"Lr9������Öw<��;��1ωI�;����\� n��h&�f@�Tr6x�쁽���{9x����u�c�d_RPn�v�J���1 2�v[��t:7Q���v�	l4��������"E�)汘[$�nkRv7��wI��6j�?졿�,�~� H�,	X6@����^$i��������r����\S��p��
�`{n�CY?���v6��v�c��C>��mT�w��3����kVX��xEc6$�K�:Ѫ	�W�kW�޿��_���gU����j2%a���k��HB����'����&FQK�v�G�[_��L�$Wڬ̆ P�&%�D��M��Y��)�|�l��ne��o|W��>����[���#s���G�drp������}�d1��0
[���*걣f�qy���寝�B	����(g�ل����L��@�d���]M����_�ŏ�nm$�M1�� Ұ��2��0{��W�����C���O}(�Wo������2Ӏ��C����z�J�".�G�{�s-�R`x6�z�Y?���#?�/>V,�ׯ]�����VL���rU��y�4a�=��=FH�k+'^�����^�l:���1[�V�>6hpI�	I��(	�,D��9�扙��O����O�@\`��5�u����ZBg=�ڜ�gfӥQ�u�)N��|�����?��/���r|�O�2��������I�.����v�ګ'�����;��3yZI�Fcʹ:�H��h7�|�JCRF/N=p���Ӻm��#�-�����m�ә&��h�]�x�cY\�ƨ7w����ɉ�_��_��~h�,c��h�+����,�&�(����K����(�����������v�iWw��<�y�" ��V��"=�$L���ȰK�L��>����	\����',#6vejqt��_�{���=�(�r�<K����5��P S�bNh8>��*�/B^Ig����d�Њ��V�� H�g��3�zLВ �p�y��'�NdXX_��{�aF��/z߿z�z�;w$�ި?����vp!��f2�G���V�g/|��n�'A�Ӟ��h� `b}$b�ʐ>.�L0q�M\�N4�="�@��_8�Q���\@k{t�B�5k�B�V�r�Ș�|x$�^I��� �Ol|l�V�]��Bk�p\x�W/ĸ\-� ��{�F�t�+��m�qw�TO��Y�ҕx�� ��$��P��5{��:6>��d�m����ɟ����������М$'Y�wLSSӂ�r%�	{;�.��X_�k��#%�`�[;���]�#��5Ĥ�E� :�s��:��z]�D*k;A�re��dt{��,�5Yy`�ܡ����Z)�EVTHև=�ն�gl9�����o��g���茩N,��ׯ����E(��)��>!b���z4!�/JKY�WQI�	�����?>�@	�(7���F���:8������l q�hSd�'|�j�r�{����u���L:X�s�$�/�����|�u�h�i�Fd$4U�4���QS�X��#G�K%�q�pU�l�Dtaf�Iq<q��i`)���r�M߹)�18�����0D܌~��uw̠��3&oy�נk	�P����9����)��;�뺝V�Q��ИNK�9a�tMd=�b��ez��*�$�*iBCAF����!�Z*;N���qGx)s%�����A7����ёC�jQ��"�����AF��q=�_!�e��v�b������u��@�0�h����e�9\��
�1/�
���6���ĲL��3��Vt�@��y.�IE�z5MMLNN�Z����	]~ع�����}�*���DV�����'g'���V8"�8H��������ĉ�s�;��}��˔�V�zW��N���.�D��,j��)n՘����]4�0�g�L ����SO=�?71;��ꉤ̱�n-�K�8�I�7�)_����ስXY��η[]E���f�$]���1.��]^$��!�c������4i�ȳ��/���=�i���J��l���u�J'r�\n��� +KJ�r^HG�p�7�nȺ(y׃c�G�3�Me�3[>�O����?�s��쳏��Mٱ��\��+`DY�yUF�qEW��l:7��&'�������g*�|�?&�	�cH`aJ�E����!2ӏ��D~�c4�cS���M�1�K1�dT�C_<�մ��q��'�L�n�����vX����	Y���1	��HF�8�36���ʲߞ����2(��/1Ndvd!�Mk��j��5^L�=�a�~��r�&'���]����zq��`Е�V2s,�V������|��ϕ�F|���@D�q�Y'�o�N$�Db��`�q�STս�0��v�h��Z���1��
���8L�_��F�8x����#�����QǤ��%���hZ&��阶����ځ�2o�v��@I(��\E�}P$-�I�M��V�.�9�(����{_�����Z۾o|"��B��ɯׁx� �P��X��aY7jG�R}Dl^#�.���#`�=�
F��)5��t���f�z�l_�A�;n��Oǎ�PZ,�6���
G(�pD�9"	}�1"�,�ER��'B�����zb���P8�φwH�ĳڠ�H<c�}������@VW։e�����X�K�<���S���q.f&�耪rQ,wѣ�bĽ�*@2�i��7h���͏����Oʲ��������6�]�U\�t~e����p*�B*�yl���M(�ss���l�`{vL<���kVw�Ȥ����y&�+*Ϫ�$��.V[˲.��d:
װY^�U�#a�,�
z�k���G�><>7�SW`����U�mW*���F�]����S�>�X-�k����PǞ~��Z�Ђ�呪+�c���?��KK����PFk�H�@uҨxuΡ�0>�Ra�nѠ`h�;%�W��jqȄ��̙&�h_+2"¾������ҙ��I,�g�]�E �^��� 
������5D�7���-+qnU�}o#���B�#��#���`G��H�1��r�m�i��B�\�B��j��5]�=�g�1���9t���0j��o�.s�|.��HBG5� q� N�������5	�2��u�{��L"�͙�I?[�B��Sx� �`��30��H0�r� �Zl�N�F��v{=�4,�D�H��dU�,��4�$��ƕ��1D0';;;輴�����(.7��;���z�~t
�~��?�><�3� �(����6�	m�c-�{��h&�SMz���?G*��b�\��+o^���b����O4lJ�:�8��er��	,ލSX^s��G�=|�)U���TR舼��KY���'��GR�*"�l[��H���'Ͼ��[���4�i�*x�KH���t=�^�v@c�~�s��ܡ?�T��^Ұ�]UI�)M��(��d�)8$	E�`]��ݮe./���6��!�Ψ�Ѝ5�$��p[�T=����%S��x�!Z���J��N(�!Z.~Ӱ�r&0�흦e�p��(�N �O���z!,^�<pD�D��Ę�"b���tn����<����&f�d80]�	)(ik�N]x��n�֒Z�nֺ��**Q��o�L�F^�!��>����J������hԋ�F��,�>Y�gy���e6k�/}�+o�y� ȶ�q"#+㹜�M��{�p�����Eyrv�Pf	FAK!=d 	Q�t����֊;TR�����F���N8wQ� gԇ�Dt�@@���tr����Dyl��P�pk�|�3��h�����
g5Z<q�;����n�eY��T��P{/�]{��	7nt[DJ��<�u��S��6�w*to�+��?쳆�A �E�mV뎋M&��x˄7��!T���w&$,�ۢ2�� ���4 �i�q����;�^�$�v�ƹn@��X����\t�q#��a0�2�&KZ��2��BK�?�5q�ީ��E�K�Ld���i���]t�9b���(�S#�����G���:�Pq�p��^#���M'aG�5���r	mLᅴ�hPAn���>�
��L��E���HC�c���fD���������p>�PE�ۦ�(�i�3�W6^=�����'?�S��S׶<��P�@,���_f"[K�
�bh!P�k�xt��z��#شS���M	6��R��N��I��w�42a١�H�!Ww:���rxba� f�2��t(��8^@�>���I�������X���t��#��I�RG��h*�6ͮBd���RKMx�$)m����X`�rT0#�f�o���ӆ%%�UR��P��6�����\'�
Z�G�Ő2�A�sC®�r=��|6�(��4�Nx(�-���Je�h��{���
t��W\+��ɱ�����} Jʪ�@�0n��t�q�8��l�����c��˺$�$��ֵ�F�����U7�n��"�+S%`���R=����>P�M�I���ܠ��*|�?��ݞ����_H�dPőhp�ġH&0�!b��z
��ρ�n�*qx����Q`b&6UIIh�����<��.<�0�HIdȵZuqq��ٳ;�-���>�y�Ra�{��1����N��@l��Jlwc<I�� i"6����d;D�����(�����A܀��P�ë����׾^ky����R<��!��^��kX��%��f���;X�U��d��Z=>�eA�4-��}�bB�����U�V��;�� .ظ����^
\R;�	1p�]���c5��
��|�/��dػEw���> q���Kp|#�$�vuU�C}w{��>���+D@��ŉ���9`c,�NiA�Ø./���J����	�Thq���|���ȓN-!rx�&�|.�0���Ņer/���>�g�$���s��?���͋�y�@1�i��Ut���+��Y��`G� �����7>�ŵ�˪"E.� �F�p���2N��I�m�Dԛ�9뇜�M=��ê�f��cY� �(�1��P�[���47�^:�&��\`6l�X�IR��p�BȌZĄSa�HM��.�R"<���`;V��.)���u� �r=�#޵���+n�V�w&��om�K���4��C���Qrl׬w�����0lؗXN�!ᐺ\&��DY���]X����j[����y�
"�`g[U
�EBw���-�0���dw*�����Ġȍ�j�����]'yD���{c�>��)��=��6�v�[A���=���C�u���ro[	E,�N!��>������{��2!����A1���7`#�sj��"����	��Μ9���/��Ǭ�"Ҕ��d
�P�D�w4%�븠8�
p�>ZFER���\�HO���1L)_�%x1P��r��yIE�&M�_�~z����r���efl�O>q��o�:���=��Ob}(���c�i�t���󣑪&�m	���!�++*��Q�x����C#���N*!�&o�����=~dz����c1/�
EA�����0�E�EX���.��9�k�u�b{����� RH6+ ~��?�����}��'%�#]"Y́�/AE�I����n�d�{������W��KIM��T]d]��/��Ⱦk܆�uMp�Uw�����&�q���&v���N�[u����]��L)�B��a��V�R^O�x.$�.��1�K��f���o.��vӶ��[��,�ȥ�©��}�t^�xlsX4�e�إ�Ѩ��i��,
�n�R��q0e�d∡*�~��\l�eM}��i�x@��+a=��d��E4�hY�m��v�L*M;�8�{�E6Wѵ��W���O��'R��Jn���zT]��5V�V��Z��H�Y|W�[�*�N��M����C?j���U��YLk�)����a!���w��D:+	qtJ�q`m/Lބl���ɰ8���h�a�70!�[��P6�, L�r7|��d��=�E�7�b�E{1�8��0Ck{Hq=-!�Ng�������s����d"��Dh
���Y*�?��NT��t
����H���0O 5I p��T���%1@_�n�Q	})G�ڴ�*�˻)����A��MDU��&\�T/����]�j	@<��󬨄Q��l��]X8�����|E�����{�s�p9�K�Z���;�(�h������������|艧88���@��e�_�>�;�V6�+W���淖.�=�o�c��X!������XE2}���!���f�/bIY$���� ���G�e- XA8���<v�[�k��X_����&w�k����vJ��:��ы�w� �`��dFFFTU�e��_�$G���h��Qc����b��'g��Txfhm�j�,x����@�j�>c`��Ϝ9�Ji�l��l�
��Đ���.610m�0Tk�?��Ͼ��&�GXF�T�g�K]�H�����z4��p`�޳����;����O�<ӗ�n�����}���Gq��M &@ٿ%.��z�$��Td�Ro��ո��[_��a�~�`����F��;����볶~]{$�>��~<e����f�	��|8֢"c$���	��({>FT��v� ���R����9� U_M����f@�!�3h�框;�#IJ� 9/�Qz�ȃ�����v6��N������J}�JI 
��
\�"(3����?2{�o���)}�c�b��j.�\Y^X�;�a�V�He�*`ǆ�P �N������ju{j"��#�勥f��b;>�֛��O�?|@�/F�16�)�;dH�*���e f��������A[�X9&�Z�^JҤ�;�c���'?�ۿ�����&	oI�N�i�j�
1S LŦ��Fc�c�E��i�\:�&�?h������(��r�Rx�0Qŋ�V�-Q���_���3{�7}EPb]@3��*��O
8�haa���ǏȮ��MZe�ԟLڿ'��N�[{�~@��bz\�u�Gq�Ng		�� �=�j!�ԛ�ڰZ��$>9��������ƅv{qqq�R?���|	Ȃ("r�T>�U�0��Z�zR���,����J՚��1ٷW���j�����?-ǎ�3��^5�M�6A�X�:#�l,._�b��ڬ,ʰ����-�W�������fr�z�nl�o����ljJ���VN �� �a���Ö'���"��9�"1���#~?��]��������=K^Թ]������MM�wmǕ��4��Hs3��1�W�e`A��ℨ��%2,�+t'�hTF4��E]|_�.DN$F� ������,��$x�]x�eK�#��h��Î���]�t捗�;<R�/v����
��� nH�(�����8�Qpxl|ȃ��S�4,`��2U5��m�v�S�d���#/����؅]J�_T0���L�-;�9�9@���1�t�a�Zc7�Np�M$�a��X:C���q2��������\[C�~$�"�I*U|&/&)��Cie|AD;��Ce��Jm;�TUI������cǎ���	8p��������t�ѕ���ƕ��O|��<������fvM>��e�V��Aݐ�xɢ4mdl[���Q,�R��b��>Vz`����b �~���E]�AR��a9�S%�V�$e�p�����[~��"iAyQ����#����
�C_A�ؔQ��w=�㔐����;� {�� i#�l_�;B�8���8���T�v������/�§�
d�<o 4EY���}�����֗���.�����J$p��9سNZ6X�T�h{�Aշ��@��ݙ ��Jh�D�ړ�
 ��^a�W���n����Y��@Ox�wao���x�wBH�En�QLoz��������a��V�IR�!��T*�8�� �Z(#l�|���V��`+�mS��F�nPq-��7*T�~Q!L�G�lE�
���Ȁt|Ƙ���m�WÎ��occw��m���Gw���by~���S�]|���.�_��?���,�f�5�_|qg{6[�hX�'�F�D=Љ7l)DHZ��#��K���_�R6�C��FN��_��?��?�d� ���s��[YCSC�9�g+�̾@%�Ɍ�2��-�C7���obX�A$�X0d�����}�$lta��'�J��.�KP�*<M�>j0����D�@�0��2�d�n8+a[�o�� �7-M�(ъC�T�~w�N$�g�K�����C�k�ZD��=����6q޽V��}E�M:�����s���TXJ
8P��	���sܐ�Zr"�i�#z�acoz!JVϠ�L�YgffL�Z����S�����s>�����|�ĔI"ia�2�dVӱ�Ѷa����P�B6Wݩ����D`��:99=�i!%3���҅J�"j����P8��v�����I���Q�oX��z�Ѩ*��l�^y�ԉ�W|`�?�g���G�Z @���TI��2��m��&!U� �XX
H����I��;#��0��㯿=��V�A�<JWq<t�7�3'�a�B�͊(	�U���M���� �.^�r}eYU ��"�a� ��x��.?��q��-X�ח�_�B�8�%ۃJ4�p�wD��J:�	:�����2�����]�����_l,ƾJ�h1!&30�����%�(�<p� BvNn;����b���aO0O�I�0�^ؘ��+�V����w $EMA��D{�>`h�,8�ϝ����q��J��@d�a�9	���u\GVQg^�����Y3�_<Ä�&��
im�z�k��@"F�s98?L��o�T.�x�/|�߾r��������{���/�q���n		�<��}�~��WO~kwc�u(I�y�{Dˢ�2���eJ��$���ޮ]�rVOi������؇``�
豒@��`�gL?ܮ5�vk��M�#�vz'ȝo�U��@��N��ե�z�4����"CZ�p�a�!����*��:���p����o���dB�Z@�"*�����~47=392��/}���K�;�s�}������_�|�����%���_���u����P�о��"��� .s�������h/ ��~$�Fr����;�ٻ��[��jhj��=����=����ߎ��p�䊢ۤ���T��7�%Aen��nu�Gj-\�����E���w�R�J�(i��<��%��AGQ�b�tx<?�~B��s�F�c��`}G� ��ضa)���}^��f'�<_Kd���PΚ��KA�>����-�T���˒�~�����O��b���i�ӝ���Ծ&cѦH��(��n�0���w�����V>��Ͼ��k@� Z�����ŵ-����~�P,�a��/��Zۙ��*������	&zߒB�pR�*%LAg&�!,M����V0��~�Y�V�A��h��nvn;���ɱN0���J������K�L{�Z�f<������s�٨�y9Ҳ� ���p/0�����6p��E7I&�'Dhpˊ��`꽨���V�{������,�C����%1	f:ݞa�,>��%�9�x����ryD��n�������Q���D�4���vd���脡9:�NpL�� Bz�4�`K-@�}g�0�������3{��X/�r4��%axx} B�fhj��)L3ciV�	���� <{��w^{}eymq�r���ٟ�x�8�Fn��*�T����5慌at�=�r��������8�?�������hL2Ӷ�.�IE��Op�m�� Q��<׳a�[�3T*�|��ko�>������+�	1O۽iW�c/҉}Vd���)p����x��%���SzId^�Uű(f����m���s��%7�~�)�[�����DD�T",[BZ�E!0! �G�+SL'S�\0= n�C�n��H�� +�+*�?#��*���6�@��+gO~��׶L��xNp=3�<��qo
1ĳ��BId��^]���/Nd�y-��. /I+2  �M����l�W6�vKC�\��[�{�,�y݉�:����@" I1�*�Zi��-�wW���W�*����Ur�.��\�JZ�kY��e�$�� �� 1��`�ӛ7�r�|s�9��s_��7o3� ��_����;�w��7x8t�R�]��Hl�RO�-�,���| ��]o��XZ�k3���4��xC��֜����RM�W��a��1�LSفB�n(*�����5�.�Ę� Pƙ���X��*�B�*@K��\�8}rne�Ǟx�#frr���.eq�����GsA�2�kӗ���b2����P�MU��J=�D$}J�$=��q�܅�W�ٕc���i(�Xi
0���}a	ym��H���ʭ)rJ���z+��d���`-�^F���\�R��~�p�_��ߨ�>��/��_k4Z�b<�Ņ���NM�����>�MӨ6[���̵s*���$���}�'�%�!^�I`��R�,�%v:��� ���S(���t�Rt�� �^%g=�Q����m�=��O�_���+��Ӿ^���>�tN���:��
�0n\�T&a�$��p;|`phd~~�լǚ�z����k�?:��^'��Ί�:�#m�k{F�A�u�-s�	�+�������.��,�V_?rltס�;��y���
z��=hDB^\Z���-*��Gneye�������ၹ�9��ԆF��7p��ڂ��l���t&������ݻ�v�<q�\	�0yquq��}���W��c�<�la��+勅�/�={vdk��%�T�������]���R)�	��?���S�k���`�H�� ������#&��Ĥ��y�M�}ƨ>��Ɗ�v`D苠o\�J�1\G��%�P@�c�C��ĨՄP��6��]��ϙt�K��d���p������`|��&�m?���]N�$�=�4}1Uí��*�3�(�l�n�DNU��щt6�0|�0B��µ7��%�|
�N)�+���b����L:��.�p`h���:�z�y6 ��S��}BH�K���"G���ϣ�-��¢ ?d̋p
m�C� �p���fsV�����r��xVX]�Ν6�]��,e
�b)U��vZ(r�����K��Օ�Ç�
�={�Zn��ʈ��>��(��
"��`8����l/�m��p��{	�(�q�%[�a�O8L?$�UVXme�V�p� �>���,  `�4&e�2����N��x�Jka��gx��W��-�{iǄ�X�CՋi�gb�g����d�/ɧ��3��>06��-+(B��(t�fJS���׾�����?��_.�7ο��Z0�%_u"���,��x2�������|I��Npm���ǎ��}� �����t��3�T����	E�3u۶�F��v�x�ѽ'.�Ͷ8��=�wa��a�$ƶ�ha0D'	�cۚ$sfkv��׿�����?�����6T��)ɖ"emK�\+��,8�������o���/|���t��(������)ੋ��B��t�'�<��k�& 5y�c?����@�e.W��ɜ�FM˄�eJ������X�����X2���f��k�t6/+�e�d��qB�-xZ�,�����n୍�,-_9rri~mq�>2�=�������"qת��N=���Ҳ,�����Ȏ	���!�ҙ.��pQ�!6�<��l�K��a�;}A�C��JL��ґo	��:8�K[oX��g��}�G�����^�~������t>��R���N����m�ˡ���@�3�G^;|�w'^�֮���׫Ձ����lם�6255���ٙ�Mݻk��Q�:�� 1�ǒZ̃���{����~����S�ʱ܀��܆D�_O�p�k��x����ټ��$�o��%�g��l�'�/0��I�%s��S�fceT�Z�)	�,F-���J,�I�yB>��A��t�~����ֳa�-S����I���x������Lytw`ɑ�_�޴g��
�����s��7���^z�TW�ܹ3�l�����i�>��/r�X�TVVʃ��w�����1������rlMe���=J�u��Rìb|��"1T�|�ܿ��;88�W���Bwk�pi���ʱ7O���T.�M��}X[Y9���_�G?�t�� �������\���Ge~���O����Ux�44QJ��^��H����q� V����R������ ��#�uVK"V
о1 ��NS��0�`��8م0��g'O0�z��!$� �דzt	���zI�����3��M�����I)'�)0 -��;�O؋�^n7ɋ�X�χN`8��}{���Ș�J���9�����C���g�ތ�1����T�A��;b��f�V�j7,L��$��  ����+� &� �G�����58ϡ���{���0Z��|�R�E%�΀�EBR�d�YP8��O(�n:T#�����[��L*S��ڙ�2>>:04�9�@�Z\�e��R�dJ��\.�K�͐��cZ{wM��g���HyyuidLCEdYI�2�y�#ִ�p�x�
r�c�P����%�2��i��� ���1[��R�4��!M�pV��,�*���\楗~ �y쑟�����Ə�c����sX�Ň	���"�($�{BFˤRZ��G�^]�?����{\KI��B*���e�~F���G�925�WS��(rJO�xnv�����G�W�E��.&�ĕ��o���3�uN�Lwʱ0��%����eC�,�Kʰ�K�Ã�������8��,���
`�5R`���R�<\8w�|��������R)�pܦ	0Gh����
�0�������;��N�����*���t���Kj��מ�0�\�u=K�}�3�L9��j�嶩)��זӲ�m�'�OM�[9�+��ɺN��Hs���%�N��\�,��]������W�������}����2��\�^T$uqi��S����>ʉ�/��#�O^�eڲ���r�4QY�lL��s���k3W���O>�k".<aV$Vx߯5M]�(*WY��湗WV>��O��j��}2}�����W[�2�����M���p�����r����YݰCxT��C����o�^]�&�F��{���Ò޵��ݣ���m��r6q���蟁�����\�'F�X����DU.̫3#�}ք#͖��F�Ϋi{*�D·O���[�=[.k�P���Q��gx?��i��0R�+Uyu1�{?������������� �SRյ,>ѫo�Hװ8��|x���d"]�s�i�(�"+�s�����ӱǃ�L.ReU�
��]s�~���[o���d���X�*���!�iG	,&�-�s�� �X�[�~��g\��nԢ��A��9�1x��q�^�cK��wW�B	� %IM�D��ƒ�8m	\/�i�V����!*�� d�֮I���s������
����'�Jd��|���c�U�f3��&�Jy�M.�&\�0�Ii`�}���)�5�Z����s�F�cO?922R.���z�Q4l#8F���������9����\�V˄g�:Hj
�9Q< �Ϙ������{nfffj�v�F �`ϥ�2%��3����`���x����w�gy��,U(
gI�b�o˲����(�7]b�C�7Q�'''�\�6???5>x���g?�	 {�巚nJ�����O�>;9x����),��/R�Z<�)y�,�7 B����lhE�%,�S���TZ�|O�з#��\\Z�U �h*��ث�*�s�����IQaA,�8n�-���zh�%O^/	B�������j��v���soO����
��{cc����w\0�����+?|�̙�۶DR�H �80�d��S>d]GׁK�v��	`�<��Ǐ�5wmv��G��z]�4�(D-	�PH4B�.
r�8pu��?�MM��L���B̒���!��,|�Vr���D�&`�U�-.^����'.�{������1�jZ�	�v�����Wy�q����ժ)�N$*�<�΢/2�YPu��mS�ܱ��X����� qʺ ȧRk--�h\�8?[.�9�j�ͦ׆�ōf6��
��[�1{��ᚎ�x���d�m�s'�ZYn���?:2�j���|��k K�<8%	0 ����oۙ�f��M`Y�%-��%V`����R�X�m�W^�t����2�Ri`v�*�cp����|��F�Ru��3��M/�-�IT������X�SGټȡ�0�P*d*k�ϼ}vb;�=8�ٴeT��fahpZ���H�'���g�#?��?]x���_|1��4Lg�ͼ��L���^�{>�MJ���xE��500���Q��0���q�����S*�S(>��>R�"ˢ 11����!�������\8Β��Xc#j��{(-�7�A�"!�z��e`�3���_a�����n��B`��[��K����!���S�� 0��	<������ & �b*�����$�(�Ġء��|ެ;Kk����"׋tk�d8����cN�9<<\,a���o�:=��C�����t=GH��:�Lд{�p�u^�n��r���$J|�?61b��U�	I@�u�I0����I�->��@(�61J�'�qӖ���GW'���Z�]�]�w H��+˵����'O����×���Ï \i����ԑ�����+3�m�TaTrT�.
%Y˨��ZAd�6ջV*5�- ��Nxuu5�� ހ² Xhrb��.f�� �x�1X=RZ��$�x���-Ůk�Tn4>>���N#
AV�������q�
� �>ϡ*Ж�$q�,d�����k?���Զ]�l�\N ���̙s� ��C�4�?��_����1�w�cv7�$���.O
��[�TN�8��G>t�Uj*�=k�7��4����?~���z�v��c#C�k�jbrU`(��,��"�Cg��}��,��<�U[5�f(�p��gϯ�.�^]���(��sx�����[Z����]ǔ�IL�P	�k+�\Q�#Q�����oܷ=�A�O�s��,�TEK5��()�Z3�i�յ���ri`���p�*L3U�,������u=2�>u0��IpX�v���\c9���Ξ;s�쩳GvO�6�UX_2���l�=}jqu���Ĥe�s3���M�����˄eZ$�JpG��`y8l:����Z�i�5%tÝ��Pr��R�gd��j�*�Q�����`�T��R���-��ؽ�M��� ٧�ھ�w��x�N�m�33��n��fR�k���؁����U�]�;ҹ�$�B+Wg#% ����#7Å��i\>��r��믿t���'�|r|l�����ڵc��z���g����h�s��<���{��,��ܕkX�2A%~ͯ<�]ۮ��?�30�{���\.#��|yN�X�Q�I�-�����?��02:~��L, �+Y�����$H���cۼ#�'@J��:��Q:44��ݒ*���_<�.;i�1���*�^�Z��.��H�&�ʣ{v�'��z5�t��aZ�	����«�(9����|Y�#E�͉�H���P��j���Bc�DV���e�C�$b$^�vm�f��dF���%����uaJ��� �u�/J2`�F�!J������ű�I����y����|V�G������'%➮��(I*�[�(r	�B%��2$�ʄ�����)m8�hk~���X[Lq����;|��u��0Z6��ƨ��͢�ݜ~�C��6>�������������Wx�pK�|��+.������	�-0��5i�g��iZ�#�ɉ)���sL�5YR�l�as���Z�����R�(hii	v���g�����7��̙3�v�BjAˌUq�;�8
�g"2�au��+����a�b316r�}����amԕ;C�#��xz-ǢV4���N�i���R	���?����v�ޯ�9YJkrW������g��--�LLLJE�J� �3r�%��A�nw�)��zn�fYl��y�ȑ0�����-#_*	�7�%��0dӹ|��C=���ɷ�^��\����<��8EY�Rǯ�-N_9�.��I��)�*˕�e�<�,�h�+�-;�F4M��`]��/s��4bw�k�$!Ǽ���^��J
y��O��0X.�3j���fXF`����'+��9z����w������ey�"D@�v�7��@/�9��H��`N�>�+�9�M�f�-�5DY�Z�f���R���@v��,�;`�EMଠ�T`=,a\:�`����j5����g�fF.��4����W��
>F1��U��J��ɹ�Z3_�d�i�	�2�'�dob3B��O#hѰ��9}lh�C��S�ť�b���f�^o�EU��T�R���#�|��g�~zna�R77!0nQ^U �����eTm���'?�x_<y�m��5?�W��,��q�������	z:���#S�����ӎk�U�n>a,,._�_ٹ��O���l��hJ�Z��6�j$��p�|���={ϟ�h���O<���C����Ο~��xY	}[�(Wnbw�m��M���и.��C<77���|Z��t1=/ oLȡc{4��QN�1�<���Z�)u��g��s���;� ��"���9XN+�pY1@�e�xp�8.'�Xw�q��6������"����/��a�?��#H{�ªk�CbRˀ�SX4EFPlq�5=d���vn +��MÂ�V�kW.<���%����0���
ָT��l�1EZp&gI��ct�m����59l���_7!������D��E����E��)��lDY���性g���K
�&i�iv��0< p��$%n7��ɖ�%I nƛǎ�ڽvX��(�'���+��/� a�Ǟ>�$�NEl"W�k�$122��2LHRH����=88���l��F%��E0a����<�a[��.^�Ly��]tΌ��gl�Ud�P����mZ-�Ѩ�tmxpxǎm���C咚��'�ov�8�X  )X^�y��2Hݷoߩ�O�9{*��ۜ}�>y�\���|�B��n����B�0<:�0==M�ڙ�l�w"Ə{���7��S�d��X\\|��pvn:%�v��&�O&�7Z�i8j�u����������{�"5<a˭�U��g;��B!�} �u]U�t0G��/�S�m�e�6��Nl��Z0y���bY��hc�/̬�n��l���y�uԊA�% Q1�.��i%a+<V��( �ҙl*}��ӭV��}{y���ť��JZK�-�1�E���TF/��_9�
��=J�Y؃x$��x./p�؞$�ȏQ�T�F3z��g��F斖������V���^��Z����ى������]�t�+6	��yn=}g2��H�0>
�h/-V��<�MUr�b)��m���Ձ\)��^�5NMG ���a�M�q��r���W��zC���$�Ϩ�=/��F�9u���O棏}�iT��g±܅�eX����[bq`PQ�,������?}���?<|�� ���K�m�P�D�+��e^�������?��V�5??�0��`/X�t:�2*;v���(_�����~t�����ηY�[�4����GUMU���WW�P�OO�vkdb����#W�&�3�f�
,��3-�/��+ˁ�|�[����.W��|���pCޑS��7i�o���}��7��Fg�)�ɯ0q�Xԅ6�0wbv8��iI�`!�孖�͊�\N��J���h ��*��b�Z��*k����}�Ƀ����
�m"J,�t�r&_�,�8o��6�\��Ë�K)�whvv�V��ګ(څ�d�۾}�
��M8xG,�cWA50�a�L��k���'	|&�LRI�� ����`ݘ��������e���JZ9%:��P�E1ߺ�d���d�XB�H��A�'�R�g��"�w�w�@�^������%+$�5b����2r�g�]WN|E�������p�� ض�Y�e�oc2uF3�,5Qr���)�r+���~t5�2��._c*K��;��i���B�iK�
@�<��Q�7[F6�?��S0fff�8p �	�š<�,R:���L�p>0#�� �:��I�I�iuuujj������=���0�V+k ����
�h�����
�K(�4[�?UQ�?ܳk[��O�uI��k�mEb�wH���l��ե4=��Z�|��={������O��c5�gU�͖FjJ�mʂ\o6HS�=�B8')r2_w�Y�@���=�|�o�tUx&	_f��b'[Mf����ŵ��Tʘ�[=s�R�a//U�W��TwN�W�f����D�H�U�!��!K;� Q-����g�s?�?�Q�ul_Yz���Z�XY����)�ɩ}��b�a6�����[�+DMLI��Gؓ�0�2r��9��a�"ra��X�6�}kqu�������j]���m_�zY�ԉ�ۗ���k�<�����+5	�C?
BQ��,�
8���E�X�o	����Փ�V��ݿ��Pj|�\�6+Fe��*\iH/[�J���9^Ώ�N�ټ��?>rza�ĉ�3-�K
<���&����<��D�� ����̷��=YI�EPOgǵ��4`M��:��vķ���2�P����|�Ϳ�]0��UQx��0Y�
̑oZ�\Ǆ�L�[�������R�Y������3"G �E-A�Xoy��H|mq�����\����Q��R�Y#�t������t��=��j��sss���m��Zv-�\E*q�o�j��L�]rL��#?^Y��F��\GCfs�����_�/_O�30|��*�L�%)=�DE嫵�h��/5-/��c��:��86	�6T�B]�po���m]ӿK����!�5f�"DD
�H�R$�J�]1ux�8.�iV�& f 08TU��b�\5&�g��&J�?�o;��
��1��� ���ŹKΗ�%�7�F����x�/^l��;vl�e��ٳ�l,��F�A�|`�`5(���L�\�7/_��w�>8 !�4���9���l6W�]p�|�<Kc�VQ�<:�fK���j���"J.�b'	/���6XC&''1��B�H�I�d�bc��K4�t5۰E��/�1^�MFN�#��q�-���(�' �Tj��^���C�.��I&>1Sy��(}G��͛�	�b��3�r�;P��![:8*0���a�)�)�\�z���hQ��Q�������~۶�^x��2YlB�DՁ!�x>#�#=1UU+k͸&�EI��JϤ{�1���ѣ��>�x���� p&mc�Q� �u5_��w`Ϯ�۷O�E�)��?J��\�`�Ml�R$��t�p���* 0EM?�����q���������'�53�$�� Y��k��;d!�F �o�Mu���A���#���:�'��f&&&v���2��5MMWְŭVm��kD-w��:���G���*�צ/ϵ0� �7'��`�ɗ'��BM��Dq��y`� /�-^�y�#K��+�K�����?�}�4��$�����ʱ���:y>�x�HK��l;�XR�m��v���Z6{p[�.�LQV�ӧO���o9Vy`xdx± ��s`�'F�����V+�mۆ��_<}��gPC�����g;�
�]�| )��nZϿr���iAr"��Jh��V>�ݹ{�e֯�,p���y,������zja��(��ȾA�K`��pc���<?����n�^KeS������
/ڊȑ����s>�g�bQ��ЭI^U�xARa5B_�^������Q�"�X��;J򊮻��ꮊ��ŝ,��{�F�ǀ�,�\X�O��(����/JeZ��1���O����J�+_�&��/��<��;N`[���ad��%�%.J�TY�"��9㳦��ݼ>�g��ٳ�����\N�%I�_R5�Ac �A�\q���sEt1D�h���f�ٯl�#�{�� ����
���x��?v��}�CT�Oq��.E$�ڕ$�c�J�p�/�,�-۲l?h�,7��H5̀�3=�i�3-�9ȡ�)�F�&���vvd�#{���y��cH�i2xtS1�^xb� ǄK�S�w�uj������ރ~�爒4��a�)��ʻ,Bz�K�'	�}	}���LbI�E^�8�I��>��d�F���s$�r㈣�=J�$�o����g���H���m-��z�������~ �7l�q�u�Ӯ��Q�7��b�1�E�<zLe�ňO�'�N������B�qGJ�ʚ�ā'�^P�Y�@3��>�n�BƁ�֯=����P�l�2���RH^��� +X�����" !�����'NT*�l��w�Q`@��a��0k����
�<�`��~���\� X���{^�u@&�O��mv�I�Y8�HW.�m���?��P.�˥�$���E܆������8�&��iH� ���s9�%��������s�z�t�_A�����J,�� ��++�[�@��z�������gff:2��m��m�������_&��g+j�bZ�@�u�@��w߶m�-�4���zT�Hu���%����Ze�Q[e�&_�.�>���sg#N�N��?��.�ߵk���H��4M���?R*��3�Bf�����'��T*+p�f�N~3(
�Q�3�"�#�b�F�3���e�|��&�A��`����H��T����HUWtrjlK�L.V@����QM�\�)Iz���Vʠo�L6JC$/������<����H*�߉u�Nܽ�kQ�g6�͸�} ��X�x5��_mLS#m�So�hnRu����4��&g�_��o���>48�h"8s�tM�y �#�78b,�Ie`�D��cѱ�|����-���:�W��T#�����`)��C[�\7<"iۓJa�i��.[,e_y�������~@�n�����!#�N�2�1��+��n���uH�u�)A��ZH�l�px��ܐc�#������6f<67�.Ţ+��44ya�G!/H�6/"<���D��@�9	���?aV�Q`�D-p���֭p<үG"��G�V��ѣ�4��^��X���J�I��,���3j ���� ;F���|N��m#ŧ?�ĕ����\Y[e�P1�TA4�=S�����#�}��c�����_�b���vc��meҹ����j��\��"+�����f1̅��)�u%�-#�jXP�J�����|���ӧbJwx�Y]K�S�&d������r�[�DO�[�;Q�7`�dj����5�0�Xc�<w|r�u������x�B�\ޱ�F�ǆ�Ɩ�jW�玾u��_�ǏZ�py�9�3��<���MF�������.�p۵o�r��e���3��rb�N
�P �B�C�"�H��a���`���+���kDµ�ss�XB���%�ǋ+���p�z�r�m�A�ى�A�Z��A2~�&��m�UA��������!�K
uI+܂�y��%�Si�ٴ9�O*Kp���<Hb��>�6���p��3Y�K���yK�{�I��V�i*��}��I�33��k�$G]_�S�V_��444H�V��|�Y�Z���4:>;���j�����'''�Ţa�)}�
�P�>Y.�Ⱦ��H.#xN�(ǌ�mުN��	�"΁���T*E�-�k{&��w 瀋F!$8��H���l��K�:_�^�p�ĉ[Y�cJ ���Q\�Q��#�!J<�z�[���b���	
ƌ|}��w�ve�z�x�P�듔���yɳ'sɋ����A�3o�㫼�ǌS�9�<
��*G� P���,l @�[�0x�g�x	���b�>�S]���F�̡�7�u=����P�Cq,Q�ʣ�>��/������W��Wvːŋ<�A�Z�2m�X r�!�q�QDX�U?��S/ 왞�ư5��7��*��J�R]�1`��s)����Zv3��K��B132:�o�.�`���RX�q����?�P�e�Y�%�tQA�I>,˅��+iY☗�!�	�kHT�d���Ji
L��������#M��v�Vo�W�-\�>
�@��;��x7�л����8"��sor7�����b�;^>�M���ퟔc��L�z%Ӎ	b^KT�*�Ä��ł��ɦ��	�ثx��.4��e�,��ˌ�kgϞ{I2�� �b�&%l�)����S�G�?��3,��:�cl�����v
�˳L�H�Q �q�F��:Nޫ��1��%[�pO��;Ʈ[�f���S�X0�F������і�Xo�*��&���G��`�{���5Y�UTBपJ��0���Ko;��(~Jdh� ������@��D ��~`���C��!�t���֌��.�cr7�$S���9δL�m�z��C�C�؅|���\6�&�q���u*�$8��uF���"A�T#̬���q�? P����O�ҽg��u��%��.�q�,�l��E�
d�dDT9�ADd�#�8\Y���"��D�Q "s+3JC�p�D�+0�r D�k8L�����%p�eL�y��c~u�Xb������7����hQ����C?p�}BI�^h;~�#G<��T1�Ω�4j+B������ |�JW�&��|>_��Œe�ؗą��S��PW�z @����.�v;�T6W����Q8O��KKK0}��r��®�LFϤ).I"����(f�0TQf�?�d�d$u�qT�2RJ������T8���H!�,�MU��hVF��wDY���Jm��P�����z!J�~��m�_�������%����fG
-��$���ur�B䣭0���d(�pG�t�%#�iʰ�G[����^0�،�t��4k4ꔍ�D���ɛ4��z֚���q-E��c��s�$-G�G�㻣��q��̮�wB&%<�v�<��%]��&��w�v��t�i�$����u7��ټ�]F�'
�{Y�͑O�o��q.:.�M��=7�-d/��t��а�[ZZ�O�!�a������k�z-��1��"�{�C�mC0L�M�5��W�N������L�+�k�*}�4*�c�9m���V��
�C�=ucz���)�H);�V�ɤa�q�L���D�������3�R�d��]��]F]�*^U�@G�0G�"�B�X6=�X˜ո�(bWE�lF!xN�p�4Iu�9��ۻx�N7���;�{��Ѝ������={vɪ����];w��u��	�p6�V9��"q`x��xvﾝ����!�2��z�ިV��l�Yo��201N)�m7�TE(�n�i��X !˫�ٞ��B./a�
%��Z����`:X�t��t�X��5�����	2vg3"V U��I� �$y��XXe'���F��ak4##c���#4>1��f�9})O� ��9�R����]3����m�*M��.K��Y"��g�nah��=_D�,�+��RL1ZX��D�cjj�J�`�����*��}�k��"iy	�kZV&��o�&�۱�0�Z�����6Ԁ�!��ZZ��� 2C��U�'ѳP���V�H"��\G���P!�Q���qGSC[�MSs����Gnxo���QW��i��z���Ї�l^��k#:J�b�\����'�+����4X~Fl��e��lֲ�8��N� �$j���0p-ӵ�h#x��(�%�=�C�V���(Љ�^�
�Q@a+&�c�V���u^���x/�C �煐-�:G�s9+7p���3���	{�,C_�YS����=l�/Ż$��!��T���7��v�[��;IR~B����E��p�;pp��؈m�H01�Y�῱�A�t��i4,���]'���Ŝ��+����Z�	��1o {���w���My<�l���NV���dT���G�@pv�=�j�� �jZ�&ԁ4�ͦs��7wx`�C��-I���`���
�rf�q�����k��N��4����j��i,�i�xd�˄	5_,�N{&�-P�kxt���fDA�ڶ� e�KF���K��l6S,1UC��� �d0�\i�={��2d���z8T�E+x~h�be՜�]z��k�2��u�]-��PO�|��]i��n9��'��[o4b�B\�@�-7n��@O���@�T�=#�f\�Pd��b��ѯ(q���`H|̨~�F<��hQȈ�� k����0����C�
����L�PM��\�L����nE,����ۻ��I�d��-z#��A�M��O)�����1���cn�6�=���!ɮF�{X�C�%D�k�!e�9*��Wc�¤ Qr ��J�`�f��Z��j5��*�<��aX�ê�����' 0 ���a� ��x�k�v������aՠ��1��&�Y�W��᰼���0�ǅ��n,��H�z��Y@�2��Yn�(���؈��@�ߝQS��O0>�e����q�f�c�+1U�F�z�}�Q�p��`���;��/���O?�y�y�g�n!���!��2�_�6֖�}��糥�G_����}���`�%�޶I�\�`f�[-��_�!����zs�Ә���m0��ժ��׷,Ƕs��M�a��?�Y������}^O�La��7kUϱ�������o�^�.0��1�hz^ ���
�˶��b�&���H��D��;y�����X�� �a'`�(*&WۥP-�k#dyyu����J5_*�Z���F��i��C#�w���3����[o�e�^t�M��>`=Bq���n �y�������uX����;��obӪ���N���k=����q��̴�,{��Z�*��J�]��]�}"�d׵�N5��D���Ѻl���z&��<`q���Ø�g+�~W1�-?���"Y�.~�M �V$��w�b�w���$u���1낵�긞P����
�
 �l���%�RbPW����JmBc����4TU/ ��v;��>���}AX�-�I����6M���ǜt9�_io�a�D]u#P���5G:V㣆(z�u����b�\�uQ�������vl��_X��A����S��YH�'�0s������E-{�~Uw�
�YG(�83�#�jJ�'���zΎ��~��]���!�õas|,�cW��o�m�w%E�$��]{�:�:su�e�ԓ&	��_���۶�v�k�����Y�`#�c�Ν��r�T,��q��/��ՕJ�ȑS�.��9ϋYk6bW��VVז����/��_��y���A����`.���8U͢�.��{���$|�l��]ApE�(1�}_�S>C�0iC�B ��a%�����I�ei���/������z�~����w?���)��|�3 r��"�ƀ���i�*�F�z�{��R�� d�6�������G�7��o8!a=�hs'�,S9J��ߘ���������HI"<-V���x[ 
�2BA�k��#n����qJl� nV�$oy�ta�;Ay�d�ݳ#��3e	��[�sNb�~Y�~�n=��:��rBy+n+�q+'��X�zJm�=����DA=�$�ڶ��o�N&�S̗M^Y�������fÊ"�X,5[���1Ij�E�X��>C>����Fb2Nbf��
�/�E�E�s��Ƌ�J��}F\� ��w<+���~�畺3B|�G�*=�ԣ���������������l�$F�G��8�>|�RwP#��4�u3z-�K;�Bd����
'o��X�g��S��GkK��R�4��i�e�JA8���"�i��lbL�Xz��g��ٚ��d!�[���g"�ȁ�O��ɛ�n�2@X�pv�8#,���rj��rz��R���FRz/�?��6n@���Wk�453�ĉ�	��N�9�?���?��㏵]s"�v]�b1f?�Aɪ�h:��Ä3Sd�v�+SUI����	�8����(�Y��p\�` aY^/8��x���j�j�����ŋ���V�4�Ϝ��^.�ϟ?�Xn�<�4�vC�ޯ"{�	����4n����$h�0�6A��_$�T4 ���(������y���o������GU�T�c�,k	�XY�x���A�U�2PO\�1�/�� �x��"v�Z���,q�� �V�&
�*3�� 揂��-J����C[d���x{x.��X-3���c����^�#��t�=��c�93��R�;���������c� R��e݌������-[�a���Y���Rx���-��n����~�u~(��éҺ����V����$N�>:���f��~=��-��~�$ �*����)MR2!H ~%��p>��#K����Q4��35�j�7,6I�4
,��k�ћ��Lu�MӌՁ:�vm��5�P�˭�J:�v�i�~�ò�NA1P��T�fRd=CBA�ۂ�Br�PS+������׈�xp��mi�~6$�Y��fAF;�4���s~ %��������Oq|�7����?<������Cӭ�X�D�~�+�rt�C���T*��t�)fj���f�qqB��-y�6ў4�\/�n�nI]vO@�o���髳:�o߾�;��^4?�,I��N�aچ�9���ħ>�o�NE-
ߨ4�"��c�O9rB�t.�aXI
V�ř�.������l��S�I,,P��b��X���۳��\l+i��B<�B�V�%C q*���PL	�%��i��-��r���c���D\�����k+��|�Kg3��D��^hx�����H�����<w�ʕ�|�;�*OMM�����kZ&LU/�k�8;���+�9�fYf[�ɮ���`XNPs%��B9���\����3�P��q]�mQ���Z���Z�aZ*=tߞ������a�<{��Ջ�b�e��F6��P�\�۶~�k�{�����`�"g0�e	̆�Q��EI��u��
�8�������v��%��Nw&0*�`�5Z��Gm;��k+����dh�� �m�n�+`]�j7�83�a�h�9�gc��T��|��R$�r�h�`J�s9���
�y��Ȁ�\��I�g��v*�^�����mn��'�����	�̰1�Ĩ)">6ʛ�1��F��@�ه�Nޣ�����.�.�O��Փ��Pas�L�F]ş���Ɋ�T�c�v���eQ~�j�(�v����vb;�Q�ʑ�&P���m�ڻj;�hM(�o96�M�a��Kv�Ȓ&���D���p'Ŕ������[(���F��ɤvn�v��qӱ� l���X�,�|F@`d���D�RO9�3��2L� cI�	�5�W/%���$�v��N9�F�q��ڜg�(.;�"���>v��[����	Q�V�|�T*�5T�Y�����>���T~���.A׳-�{�����g���}�Z�����|7؈+�^.a���������N n�nS:=^����Lr�����V��z���<X��Wf/7ͺa�XH��AHF`�U��L��e;TZɍ����ON�ow��1��&&&�m�'��!챒r1=_"���&8V�L��W"(�Oߏ�t!b��-�j�U��*�����B�j��ұ�ZZZz��W_~�o�y�Qo�w���_����qiz�?����g��J����a.D��i���a��b]2'*��)2&	�P{�f�CU�6�7J��ܳ�bf��h��q�]=x�-��F��2�C	PI#A�Ri�6�cRD�sQNUD�u����o(�s$
 v�����h���*�mzC}��t"�C�1.,�+3��E������v�?�((�5t�PW�lW�D��R5�Z$�X=L�,q�:4��%^�r8�xnv��)[���EɌ�R9ܭ\x?�-�㛬쥼PL��4%�r��vLW{R&%�э��RC�����6
#b1Q�>�	x���Blm	�B9@V���"��)
`-M����7�>R�}�߯t<&Y?̄>�C�Y�"q�R� ^�Шq�BqddHK���s*��bӨ�����8	i^c�;p�����.�V����C`OT{�#���|?Vn��j{dr�3'=���B�x'�c�O�B�8��EQ4p\�m���ւPq�DނQ#N���W>�K���?��r��E��s��y�k_�Ə��K.FC�,��<���m\���N���ٻ[�:=�w�H�-��4%��e�L����5�T)�˳�D���g>�Z���k�B6_[������2��=]���������ghh 'Lp8����̥�Y�&-� ��T��2�|^�Y�,��ҩ�A$��n��� ���b�@H�`��-� �ʏ�F����i�$&��Z��ڵko�q�	���COO��Ʋ��?�0���=�\��ʪE :j�ەzρPr<}�B�D%I ��V���=�H�Qʍ�	��wX�W;���!&]�L1��g���_�D+w#I���R�7G�Ֆi��P'�#SW�+0���-�hY�Z8��2@&8yح
��xdA���:5C�:O�*8�����jЦ����$
�p����^�~_��9���\����s�
A#z���=��'hc��v=�Ou��aN�]j˷	��j:H�M�|�_�=�Vp�P�|�8�Ϻ=&���i�m�̍���CP >9MVnӔdI���)�Y���0�b�H�Q��n�]�����)�`155Ų[��I�
v�G��A�(c[Ww���' F�|�R[�z��uk&3���V��`죶�V�TPJT�k���xUX"�Ixݮ˄V3)�B�{�h������Ν���fuQ�k�<#� �TE��8�1�y������ӳ&(K�-��U,&:�:=�4$`����i֘� \*@���.�Aw%�jrd��յe xcC�ݻ�����#���/~)[�m?�%?�-̽��W��_�W�S�><P���lUձ<���C�"K�~T�E�r��7)��{mqOL;�N��.mk:s��p�b9������EI�uAQS���J���?���~�SFc`HyhtvfF\�P�
�zeii!������ә,N�n/^����7
ebb�)�:�w���b֫���t@��Q2��'�|lKR�(�D9/�l���� �����|~jj��l�d�Ck����QYV'�'�V�1�P=�dmrr��O|�G������NgC�c2���5��e�P��ׇ���\P��nE�]�#��c)M�5�u`��"I�,�Z[����,/��WWtR�aKUH	�(����0"���=�ubbR�1�j�:yvv�����}����'>��m��Z%�J��pn���5�:�2ER���G,����p �lE̟�M�>�~���L&e����.��5Y��]x���IP��,Dd�,�v�rn�Gg�.�3���5�:�?��)O��~�a H �X���֯	�����JB���a��q��p��2���c�[��7;���m�����K<c!�e���{�����J$n�.��_/���O��� j6��F���]����S=\��a�`��P/���*xN+�/�
|��CB�믌(�T�b@,q��p����uY$����R{�u�͠�\��'��o�Qx��6�T�ET���⸚����\�r��S�%3:���ѱ�\&E�X��&g�Y���<�����2��Gyx�]�N����}�;���aX�,F�ٱ/�
�2��M p�:�Hd J�
�dy�Ķ��Cp��+X�ԩ��Ɲ�h���b�L�8 �0O<�h6��|� r����~�K������m;��Bފ�n�(�`��^y�?���u��4GFGxpc"�LU�9xl-��o����m��;>ʶ�B������(������6�$��N�u|-��8B��g���'0����z�w�o��sc�}��є*�799�s��mJZjpp�Q��@F�Q��P�G���}A������Bwp\8�
��ȝ��F5r,����o��a�p<��𬡈� ��Wk0T�bDЎ�]JI�MȘAbu��e�ZƐ��V�v(x�l���B�l����N��r��K t/
CU� WH,*���_��_��O>�Y�0e�Ŵ�Ik��!��(��P�m�*(�*p��5�:r���J��x��BNݫ������]�f,޾�h���O<���������Y]Y*�ʼ(����&�E�o������\.�
�>)�D,�4�b]ƈ/ M�� �d)�daem!�B>������?���ț�-��GA(��@���vK~��rojՈ-h���T�G/� P�xtJ����F���̥��twyQ���>�� J�mH��s��>�*�oW�F���p=e	�U7o�I7�,�D�E��LK���&��PJ\@E=?��P����A�8�N^���zn��v</&��ϗ�{��{УZac�R����'�b��k�hSsD�F�C��	�A�6j�痀N�dQ+U�|ֈ��HV�F��+�4�|�F��0N$�����ϧ�8�HU,��Y��u����v0�d�B�'f����gK�����߭��<A�4-ZY57W�]y
�¯p,�I�8n�YF�8�p��6��	� ʇ�~�<clx�(�j��z��`]�$�b(-����y���o~�����?�n��te����1Mozz��_��w��xV���6=Ǖ��(!p��k�|�\�":Ic���ڏ4(Nt�b��a��$Վ�"�;	Yv�0�I��"^�f��g:���-���?�.�����ݽg����QDp�R��k���ס'�SԂ&U����!�X$)YD�����������Ͳ6����,⺡i��e+&`S��"`E�#F����4�5��E@�i\m4��!��?�({��3Q�@N�0����_���:;׬��<z4�)�Z���D�#���q�-k\r���~	9aME�q�GF�g�_��o��UF�b�&I!AN�Y �klPg&Ϸb����kD��Hb!���qV�806:?62���Lӑ��������/}�O*�5�ϡζ�2C�U�W9!��~$��r��!��~I�6������,�_��8����'?�I�X�����<��>'2�F�E��{L
�Ɣ�Y�.�Ƅ���$��.*�c�5�r��Mhb�{��o{����jM���
[HQE��W�����I]X(zoo�d�3;���Z�R&�$)�;Ǳj\�g����O��e]���%���F$�~	��|�e7�+�?�(f�#�1Ie���b�6c�h#�wl�ct�����-1`��Q2#b�n�Ն!�q�bOֲ(%L�	�s>� �H X9����2��͋jq�Ȏ��V3�P:O�|T
�-�2��B�Ղ���O<����G�i���b�ut7��OO�~ɴ]����K"g�rv�����u�-����+�"�������mj�_�Ư~�~�S�篫ٲ�y����K���w~��xقXYYE�?^`5Ad���ͧF�~)��N�,��;y P�t�.��l�M�a��ಈ��28�b�կ}�왋?��SO?)Hb�����dDvn_EU1�xA>�^(a��ɷ�F�VC%�j�)��t&��Qg=b
vP�!����&��p�cc���###�O�!�Нc��˗�)U�?e�Y�BB�B�@���)�Иk�CUK	�b��*���ڹs��<z�Z�ÌJ�R���j�hlߡ(�{��0~LZ��v�-A;w��Ѓ)-s3ў�4���G�c�l�N��G���Qp�v4Ϫ&�l�#+b���O�8�>s�c�'��@q@�`!C]m�t�bq�#=
�����~u�j�i�Ɗi-%IpH#�W����zhFW��,��``�������E�])M'�OXz���gSH� ic#�g����>��On����_��|N�e���=���P%3?=�Ȼf�Α!Z�]X�SH��"m�G0	��6"�.�q��=m�9��q����-ǋ����3EaW+�]#���I�T.�+�Q��\:bӦ��N�t*�/0����&����,�2D|:���@��{��qQ0�
�`g��c.)� �t]e��dB�M�%D����5��+'�YGA�߮]m���_���&�u�B	cxH�-0�4��}��F��Ƨ&EY�C$�!sezưl���<�b��gEi:/p��&J����D.�q�`ff��_�����b�-Y�E����V�8��q�}���m`q2��w�"ߣ�HlB4PP���/���}�]e�������[2齐� �	�t�"��"kY˺����U~��+�� 芀 ��� �@�$��L2���vz�����=��IBB���{�q���{�w��}��-�{�q�W.9���LÍ%7x�խ?��7֭[�}�vJx�"�#�O� |-Q�;��I��ƨ,��3���TQ���kћS����"UU�v6��p^S-�:A�v传C&`�&t�گ)���ʦ������?��-Ȭ���V~��d)&#q!Y�J�x��b��q[V2�.}�.y�./-�t�@D.�}� ��TX7�Jѝ��DP��Bxr�$�	�#�0�T.�Zݲaaɥ�S	ET���Ÿ9 W�s�@9�q����+�����?QF�^ʑ�|�qߘT�aX8��g\�#.��1B�9���Ͽ�2Z;�`�|TU�`�ٶ;6�S���%�����$'R�S�Έ�<�/J��cc���ָ�J���ٶp�LIK��D"��=F�K�� HH���s[�Y�rҩ��p�/~�C�>�i�K��&^�˦1::<�?`����,Ù���knn��K�X
^
a�W�*�q��@RU��lC��EKn���!#�b�s����l<� �^%����,v�1�R��"���Mu���E�2G$�����*p��(jR7��s	M3�<ZE;`EIuT�%%�|e�!]��x�a<�?e����['8i=ߤ�>�U��gذ&��N�j�P�#?���"��v��@?8��<2T<$KR�ĝp.Si��b`����\@�l$r���&��Y�@��<j�x���ؗ�/(Ů�(pD���[K<&�����R�?�GL�$��m*�-y�m���Tf�T���wX�zh�Ԥ�*�b"�Rn�i��lF�u�Ź��V�,�Jo�
m<h�.���VR=�C�F�I͞�Ӿm' Ǒ6�ֈ)<���h�m{>���~)H �Q��h�<���B�4�,1�тJ��c4h�C��X5{�q�6/$���o���c��a{ڷC�l��p!m�ohh��h�hrtt������4���t64��S���z�I��ȀD�a�G��`�,2L:.�R�ƞ}�	7~��'�=-dEX���X3f��۶�����y<��՚�LQ�X.J�{���@�h��aE��9�9fJI�!�b��?i?��&1`�ƈ�YD8�C(�D��d`K u�9@�,�� ��i�k96��ށ�}驪��׊"��S�:$j���Z^T���8�2�O�K�2X_�a<�L&�ұ]�Ʊ�!����b�`���҅���/�2��j�1,����V����ʐ�DULp	L�+�I7�
�وФ���c��_<6��5��J���0�!���[��7>�L��$�<�B�
"c���5CG��1�$�`U,�wX
,K��s���d
vs,�^{�ٟ�����m�d5S�qmKQe϶R�����T��+�K����c�? �W}<
j�p8K�:Q�Mػ�mL���]��|#�I'p8q��eI�-G�ԳΙx�y�Λ7M�5�3'r%�P��f2K��*�je�>�7&[9����84� N�&Pu���!A������*�픍	xƂ��\'���5��h紌F�����Ś1Ǳ�M^���:�H��R�xDbo`)8��{����Y%���c�,�	��L��.#pI��(K,��J�v*����e�~��p�t�)�r�}��7�6�O 6��YQstB&��#g<R�x��IztS�;��ѕ�k�ē�jQ�j�����3W�B *
��R>��H ��;U�ᅞ֟D D����bɩ��b	
����$@௽
7��2!$��Jc��b��(y��X��Q"����_��/o�Do����xu�H�@�����!6���x]{�&u"��Xyb��"p����7�t��U�}�����j_�S�%����'?:���?��,ŀ�ٽu�C=r�}c�$���?[6���A��h�\-�?����K��d�gјr�ܩbA�<z4�A�-��h��T*ъ�#��DY8�]�4Tm��$	IRȆ�H��'�wZD-j����(z��1�ľ�%�̥q�	���@���R��"�Z �5k�"��w����^�ֱ.�G
��5�A	|�X�W5�4��@�C���)�N`���&t	��]�]0���s�����hkkk��v��TUtS��ys��s�e�ƦL<��
o�D�>��*��Y6#����#��Y"W�����	�������%8`+<��D�)������s�-m�䉪�)�E�Ƈ�(��+ʄ�����*�����c>o�/�I��1]�!�yL(���[L��e��2̄��6Q�<z}�
�2.y��>i��,ઠ�/�c�Ԙ������*,�t���?4s8Z4O`$��G}e� C�2�,
��HR+!��邳� �6�W���뇀:�~�i?��bb
A�Ӣ�G{]9�L����Kx8�\k��9&D�~� r��hgsmD��t������%BSM+��Sפ�2�f��aV�T\��|� �.�$�92}��3�y�2g4UA9�ez͓�^�p�Џ�0D9;$�M��({�O��d���	���,
T<
��x![�UU�|�\��\���=p�<�Ql]E�~�勠��5|�!L��"	�ijI�s�^�����P"U�8���*K��	gM���%�,PE�����`������x�w�a}��w�fy�1�hG*�8`��1Վ����h�шX��l6�qFM��2�2{�c��C�ߣ͏��H�U�d*��'�\�i۔����X�y��k���_��^��	���*D�m�M#�}4WNvjE��[�w��?,�~�|���4�C2<�혒ȶ����~[kk�;v��M���YY�dAH�UY�����3�p[w�h��rL90B�r�f�Z�`~wߓ�.\�K���᱂�eE��N}�aCG9���'�s�veSɦ�$������aI��i�A���`�K�l�fI/+��m�_/�w�n�ֳ{�+�瞳�:+єd<���ő�ľ�dA9z�"O:co�%q����桰/��F1�Q�D���Q���0���d��⒠�a�0rO�',�M�+M	\����	R�7�<�C�iM:_oਆ����QD�Z�����e[�� ��sףm��#,�!��H�8�,å���" z��j�JpDI��H�0굨F.�䜥4	W-O����B�٠
�L��4)t���E=��,^��j��R4�ʘT}}����hk/&�Fԛ���|�ma��!S��ٚ��/����Hcl�԰)��:d��l�(����$��d�ȸQ�d��&IDTKZH
�A@6B%#Lg۶�=��/_	<~�����C"ca�I�O�W������O�o�	�����q�Oc�a�P��K7���b�ǃ�����K\���t�D� !}�p�cˏ;�ʫ�W_�~������X�ʏf"�:�t�D��Μ="7:�1	~�u�j'P	��ʔ�k����	kE���b�CF���58����^��U__�U��V�*� ��`���A���۷o��Sv�NF����f�6#q% ��>?�Z������3,�w��eY���e�/�;n�_}�#3�:��k�����~�'�y�Tv�2M� �
l6�)��^���w�1{v�aM��Ƿ������0�\M�k������ (��;^�HS�G����J%K�0p��E�v��]{��[�x����{��رc��>8u�d[������X�9��x��3g�%SJ���z���~���_X���JW�E�ʕ��

�I`mIG�ՖP�����BR\��ƞQ6�i��K�U��d�X �����9/p���+���]�=Ɖa8�v��V��z@[��оﬤ�������~����H[��N�ڻ �XaZ���W�	��4���� ʡ�3�����be�\��eC���~�������uh3�).���k6?���z���J�L�8�"�7ϑ�ʸ�"�H�`[t��:D�������xϋ���)Å��s9�z�ZT�6I�.Rߦ*R�p�ձ=���t	������r�f���=ҏ�jJ.�R2��2�َM�I�偝�l��c'�?�����d�*	H�(n=xy�k����ӧ��dP�u۶m'R>��+�Q5=^U"FA@
�(����^{r��n".Ɏ��������ŗ_���"����gɢkfp�XU�-�1q���}1c��T2���$R�h�C{����%[��aMӨ��Q�j�ف�GGG��N�MU<)CK�������ACO�9�>-��v,�N'�	8�%@����	pGj�����Z���t[���hS9����1�.bi%�0��o�tP��?�+'�5��j�+!1��H�k��pc� ��{���/���O|��k��&t������w����ץ]o����1M�lOw�eK\��뗯Z�e�/)�z���s�����O��k��;v��w=2 A�w�,Z�B�`����;<���s>�/�9�W���'?s�9kd64
#��6��X��۷G/�_ɗ
��\NV�M��ä�Zf�lkT�Y��58�ګ�.���\�Է���8c���<���T�=k�G3 �/�qo��0,S�E�sM�LjRsVa|+�M5�Ӓդ�8��I<#�e^dl�1tƱmA��ͰQ2���`�o��m�*�?����a����8����f˖Q4��12��v\��Q��PB���ȡ��$�����a2U�:������2�ʺA�O#�`�i�������C�>6Qb��"�d2	oR,#<�fo�J���G�p����\��ա��F�k�Am�[Զ��R5���ȍNʱ�:T$�d��`j��59��쁧�n[Rd��F�F�&����.P�a�M��$d��ԎUG�id�DV�f9�T�o��/�%��w\�ȱGYG�!i�a�/)C����p�O*�i�c-o|kN�5y��zf��׺�x���N[-��/n�KDsB����T^�~UU���X�r9 � �_ڸ`���}�;w��Y8M�[��׾�|=Q~�hJ��%�p��w�D���8�u��P*�(�g2�1u]/�L�8��|Op0�@�S#��o����Km���z�sGGKzK��o,���Ʋhu1�+�ݨm����yL�㌭�wCl�p��[z����غ$i���jIJ*��Molllp�^`P�-?>��J�m��҉�k�K�M{��_ٴq���9��ͯlݾ�K����6�~��N9�.3���^���/�*mbb&�L_p���x���S.���x���ϝ9{A�l�k���ْe���ۤxZ���T�%�3�3Z[f,ܰq�Dn�Xȋ��q�����{p�����դt�������x+����^Y�z����9���b��]�VMa�[��5���1]ԽB�z���{��!%2b���0`"���p淼UWp�o�ؔz� �a�7�~ C�>�cH<;Щ�
������Jd��[��Px�L�vL��X<7Q�t��	`$r|E}��^�T��+@���K�J% `��J�ǂh=]Һ�V*�#m+�fRբ��f�ۤ�4*n6U���HC�T�9�WD���JS�M��OMM
l�F�i����&C��K��O���S��g���'��>����+2
�!��\!pc	p�l�hR].�HS�=<�B����4�6;J��B̐�"i�����[w����{��cSS������fڳ{ۄ6R`��٨�;����1pkl�2À�P�X�yp���^�Ȭm�c���m��c��N �񄆒�b��r�Q���a�"޸m�T���r_�L�8o�p/�M�J-��Q���?ajJ���ʍ���`~J��(Q��e�6&�6J�(|����x���f^��G��q�a���}d)����t����D�S;D��j'�9
"���	Wq2jg�� @8�L�\�ql�"�vX,c�|sS�밒ħ��'�t�c��ѽSK�:��f�u��x"uҩ�������N?���'���|�`��Cãw���޽����	�t^A!Y.��/��1?��N0j��!�&b�n�D�y+���ÕKfs��7�E�V��:[�����~����ޕ7tN�Z�S�F��k�oh�Y��
 Y��8�q����Mnt��5�׷G�m�x�	@��!���R�<��Ȭ��A��Ѳ��-�':;�n��{?|����q�4&��ɫ�|���yK!�J]z���w7d�e�)(b�xN��W�q��~�S�T�طc]�6Ik�.8��UE '���m���e����y!M׳ꔕ���v����Aϵ����z����FM����%*�ٰa㦒n� 0@ϿiEGP�N&{G�7}zk{{��=��cP����U�)���Ϛ����:80�s�.]�c��m�� .���T;����GG�\���G����T�U��S�h=!v����O�(���G����]��Q9�(���͟�dth������L"n����	*T�(
�x ���fNw����c�nٺ+ 2�ʦi�&!�*dTWygۯܑH�W[��׆iW��ᖭ[v��4)�T�$Ajz��.S#%�L)�T�x4O��h� ;aX&��Mݥ��FٔU�4uG�������L`)\��\4�9�(@�]*�z�rɼ"L$��c٤]���&z I�j�e�p
�0�-S}�cr�h�!:/�K��)#�T��b��y�4�7�&�������I��d:�0cu�؁�@V�CE�s��GG����V�0�6uÿ[��w"+B:�
�����M�鞐ΝE�p��Y��T��'*i.��p�ȑ�_.d]��1w�AX�"��s<\2V�P�Tv�u&�B�ؾ)ړ�g5d��$TsCO�U0�������ڸ�yQQ.4Q]����kx��3ft�XIK5lzi�Ͽf�>��h�&FRq��>�.���+أ�#�R�x�0����s���.A�V�\��Z�e`"�U2�����	u�J*�LxVa ��sC��z��ϑ<�d����g7���K���栿���~~:�.�y.��*\?Sv=�PN����ғDMQ2<���8^-˕E)�o�e8QW�Y�T�|�(��GU�U�(�����J\�*�GmUy:��#�����js����":WU|�����@ [#p��Y���(�Eꊙ}߿/��Ҁ�"?�.;u̕M�0�P__������o�V����J�Q��Od?���7<����κ����mǓ1N/�����Μ����nzy\�2��yr�HJ��ø/�Ou0�&r4�,J>¹��Q� �E	�/g�
v�K
N$x+2��~^|������X�G!8~�Ri�T�.b?�jQK-�9�����Ae�Ԫ_E��P�b�X��8*%9�=�4|K��6YN�n(�O&��3�98t�m�"���������lVV��F v���>�(�-�Z��n�e�c��Y+�qY��k�^u��h��ʍJ��/�(1���͍�g���W]��l��n"��z�k�LAPR�C`Q�|��xW�7�����r���
�w��[��c��X"mN�9�@�2��,qNb��_x����'o��Ͽ����/�;G�<T�i�,��&��m�����/~�c+��}�o��_��x.����V�k4Z���AT��r�}'p�>��:�"s*m��T�-�M�z��R!f�Y=�tB<�N0U	��E��T��r���H��Ѵط8H�E�6j�9�����"�}�N(����#�&*j�y������Z�F3/��c1��áO�ե����w]zތ��DR)ʾǥ2��z�,�Xܱ�D*΄x�D2�o���a!�w �/�����r���H�@\~@&[Tmbp��y�D�h"h�����/%ٴ��t*����uixE��Ђc[�(h�J�ⳍ��e�a��Z�P �'�v�`1�X��u��,�S�r��
DQ֟D�}�h�e���D���D�8)�)�(��@�=�_��{���o�{�䆲*3��{��9dw �g*�d�w��B�8�l�Έg�XE��F�tZ�q�����~M�(dF���z2�,��"� ��F?D����ݘ��`�l�94�H�I�l�PdѲ�j��<9'�w�Q`�-��Y�v$nm����uT�y1�Æ����T:��]=�T�-�	��/ ���� \�,	� �\�XQ4�.#x"<]X1�Y"�4L��A��@�9�4P�k�����8pLO&"�&W��ǂU*"��4�HBi�Ο��&��@xCQ�ڞ�ȱ��!%�(6@歉�j���8�F�+(9�	��C���f�ڙX>�$ ��c%/�GQ;�z�P��J7K�H�iXZ#\�f��WG�Z:,n.��à*��6���S��:�7���w��^�d!l�{��;o�#d���vE�u��i���9��W[x͢n�cX?�����o�_���vvvrna޼ys��}m���`�-Y���������.;n��ï��&m��˹��~0�Yg�]�l�(&��Y�Ǉ��_�p>X��'�I��7,O�i��-FR�XC�����{����O|�SMӦ��تW75�Q*�<�T�gȒ�x��O����޴L��/��K����o��Ȱ?��C�l�����E�!�ϓj?V/QĎ���l�E��I�yE���Bv>ΩD�@�D�Q���iIV����$�JbBLM��#v�wMPx)G���_x��W�P�P�U7l�K�/��S���]��7���P���A���:�f,����!��~������X�����J�́�+�0��.�LjË��D\�y���cVG��ϲ�2�R{�]M�}N��ls!@�`�ϣU��&�� ��L(�DڛD���Yx��F�^�|��*��V(�pW��;+X�P��+���'Qĝ��#xai~��ΐ���Q���	��m{�d�_�P������|��N|z���}��[���_ ��rɄͳv��]�ܹ����o����rV&�.[���s���\NYB;k�%]7����=�� �4�X,ϛ������.87�m�'�%�`�4�>��Sv}%%�� %E�yZ����[6�{﹟g)PL�2Xa8x�У����kYe�g���h�������tt̾���M_��?��05Б���l�gyE�CˁwZ�����n͚3R�K�c��0*�t��̓�B=�\A5�B
WJ��
���ۋ�5J�%�7#��$Љ��0Z�_�vTq	
x*O�d0�U�T��f�36ը��;6+@rV�2]��lX"���]�x�݀��UBdݘ}�|ő�e�򀮈B�\cs�q�NZ~�;`=�llĹ! h5)r18Jq�Sp"�c%���S���YѲ఺f/�������?���%,ì9��3Ź69�D�8`�a4��{���/�y��?6�/|�{?�����\�TRd����v��訪$zv�����W_{5�dǩ�VW ���A������L��a��rf:���v$Qr\O������I�H_2
�<E���1 <D�/:�V^� ��x�j@���$�pj��
�e����L�ATP
������u�'��ѻ�\������I��A��#	JZ��M-���u
�kS��&E�g& �~E�x��J8�څFI��dY���&���o�&F�R"��-$�I5�8�ձec�����p ��@i���:\D!��C�Ā�uW�ܽ � ��q�W*�
h�lb��8�H>�ٖ>��1��m-ˀo�d��~�?��<�w���d7���Hb�>
�
4!����F��l>��'�����l
�jB����X�	�|�8�w�0��b�F%pm`�oJ���������L%L�wXޣV��J)�}O�L���F(]�t-��@�@�Fp�i[e�h�Ke���S�}����ٽCRxI������x6ې��X����w����K@�Vx��u����Xq��'�|2 �p;::�M��0� ~d�D���N�h�7̲,K���8���xb[�A�ր�~�ɭ�^����'��r�=�ܓ�k˗//[�X~P�X��������YO?��'�=�[o����Fss�����zx������o�t��0.H����nAg�:HmMϡ�>L��t����K
��Q�E u�>ɹ�]s���A%���1"B���c��{,TUݕ�$��~/��!��M9(��[�.$Q��l����*�%p�TU�C�k�Fb��Q� �Xh�>��O|�k���K�%y�o~�v/���ڕ+f�#*_~��G{������K�~�ug�Z�|�}���{�(N�sHY<�б�d��c�I	�% �#�����0��ku6'���3.���l:�����v�|�w?��K�c�Rٲ�'<+Pv��^����S	�֟�ֻ�ɤ�cy��fY��[x�胬��\15%bZa>��h���O~�V�:��7�M$	%�u����k�W�đ�~�4|W$�ɴ��#	QqZ�Kp�)���.���+�M����^{u'#q���|��۬>��^sX�d�����)�(��E'����-'p|��	��s���	Ա�D��L��l���}�ʫ����Ccy�quu�K:�g2��$4��K�)k�L�ӥB��^(�����<GA�Ћ�S剪�^�8�Y�؜d*u�՗�������ː�I��8X��d�g�Banb�왟��]p!�L(��J�l"�aQ�t�+����G(kr�ԡ�ȅU�@����2���� K��qSX|tD8����h�|��� ���w� .DñU�h�9����2
��w<�nzk�ߙ�k6�v�f/`�D�lX��8nႎ�*˚����_�ˎmf2q�V��(TE*dz�j��QF���dӰ�	�K��>��K�[��>m��xA��9�˱���=͍M��F�B������ʚ��v��t ������%5ɰ���-4{8}��^���@�d#���p��������)��{?l�U��!��?xûg�[�4�eaw�>yuWg�g����=���|�.���Ӈ]Mf��3a�0�<�:�i`�$Q.�<����)�Yφ���� ���d>_<B`���H;��d\5mǶ�@T5aS���a�<]�r(� 3L�|�lY���$+��%���D	ކ�$&p�M#=��8�J�����@D4X���U"1��j,;�� DA���v�DÅʡ	�I�j�<�!nf�wI�
��(	t�V�辣�L�G�J��ZHh�#%B���+�O���M���İi�
q�30�:}>��Su�D�����4-�4m8�����d|�l���0�T+R�ǨÖ�56��cqi2e����t`AU��Q8Mu�W��V?�I�P��{�3I�;,�lQ��V^���Q�����i>�7g�U��/_������ d@�qCh���\.�8�&(
vI߱c��-[�F�GF�v����2�gH���6N g েR��ʶ���k�J�Nܐ��!��,����2��#p��X��a���K����'�x�����u��j��@�d�x���	�ջz��J��὏�{LSw�N˴�uΆ]Nϧe����{V�74-^��ƤyNN��#6j�Xr�tl۲Lsbb�Ww�����r�R���r���a��׃��u�E�P,�������`�����#��o���?<<���4{^�q8�����a�LT�O��8����XF�D	�`��L] bqt�c�EL�m����X���W�� ��}6�E����[�t\���J$��bU���Tg���{,�(�<1dP0	�7l%��9�_����i聄��=��+W~���e��9�l�����[n�WJ5Y^�n�|S:&�@qh���~�k������"*����,�44{�����'�o�����i�������*:j�k�%�-�"�u@ɘJu]{����^�W^^אd9��%��N>��g�'�?����󘽐-�֮9����l\/~���1�y�S�*��ڀ��l�ô]�6�2��5,���t��h�*O �ݺ�E��Y�ʰK�l��
p�G���&���G%a��x ��eys�u�tӍ�\vy&�fA>�J��X�P��豹"�(������H".̝��o?�0����yӑD>��q�[�%���� j���FQ_,�K�ǲn�,
e�x�M7��qx,p1O?�a��[{{�$Q��p�"k{��~g͚��sǮL"~��Ϙ^�Ɯy�����׿u�=��L�#ƼT��S Mj�}#eM:���$�.��=��9g�I��ls�s��X�Q���wE�^��c>cf��y�\{饗�뒋�P�un�k�o��W��{���aT��~C�%J��Z�=�Ó�<�_�з1#bEHQ�E�6IY8�z��-��F1�L�{"�m̟��ّȠ��G�w�e�_x�Yg�u��In}i�O>���}��x�^�;k�9g�&0������_��Ww>��S����I��Ǔ��C�*Á��@"I j��lk��ޭ�	�+%�_޹}���'����X�p�e�{z�tu�lmi޾u�ϙz�}�{��ATҶ����T���<������׭{LVc�ɮ���(���=�l���~O��q{����ܧO;s-|cKc��ŋ1��q�k�b�M��+��dzWk�\ ���8��cN]s�?��?��/=�ؓ���؂j���(�zpz��`a �,YC�
z7��[7L �,	��Ԥ�?��@�PG�r	��xA��i��W_}u��n���}��`����d�1z+�PxY�T�����-XyO�s�;e�¥�a��M[l��5M��ǆ	��{:)r�
L	�=Ж0�l/R�Å"ϊ(����;�h�)� �5s�"��Jr�㨩9L�38>�UD�r
,�8��Є�3�+�C.P���Q_��Ԫ�Cn4׋��T�$?������V�f;T S���Ű�e�������9 U]��8`1�#�~���-�.lpɨ-��;"����  u��������@�,�%�_����?��\�h�F��3������0p;
�$�M͍�8gw� °r��rJkk;Ky�n8����l�o{<O�$��`�+v���&�z{zv��Ǟ^?�/��N���L����k�v L�=B�*�<�=�T�7XӴ�D�rcÃCۻ7o|�y��0i�s]]]X��i�{a�����bJ9��پmǶ�J%K�� m���s�Ř�eî�۷�S��l �>�JU#�l����E�!a��K/n��"�������c@��Z�����9�v�&�G���t�N��`\���Bab���e�̙p[�kȼ3:20<<L�}*�<�rZ�N�=����p�CU�]�QEC�ulP�$1�M�����<
�	~
0�T�G������J��^�#��>&���� �@$0�Εw품ʯ8���.F�%X8�1�HJ	6�r��y,_X4�5<�K	7dkcdZ/W���ii�7�G��X��d�;�]M�T�i`��G��5|��;����.<��w�-������?	;�)��ʦ�<�z��'�p���Y�V�~��;��� �r��"p�H�ڶ+pf��X&��&W�\2gV��^v��k^v����٢�:�y��g�Lo��}�����_}u��$�u2Acc󻯼��}&㔯����;�w��j�y�ޤ��2sH�3�PSͱ�H���Z�Np�#��XL�I>r8q�2u`��3E s*�rB���A�ڑ2�4L�!2c�쎿���]����d�~�`��?���G4��v�Zq���V������y��s��Z,�1}��}�s����On)����3&&&���$�2N���a��E���T����5'�p��s�#.#|������a͊$���f�1yIH$bl��� �sӍ����Y�w4EZ~���<�+<�ؓ8+U��i�4�Ҵ��J%/�W��^���0<p�5W]u�꓍���Ι����[;����_Y��|r��.����\����3�R�œ�n���;~��[�0I����[���~9�N��"\F���|#�*��"NVX�0��, K��u-�%����B������q�Spw�^�=8��`/��s�l���`�Y��	�r3�����Ej,���y#�'55�J���*u��/:���O=�{��������bgǌ��<��I�zk��@h�P؎H�� �	`�<��0�Ų��Ǟ|��BL{�O>� �e%z@t�Yq�ٱ��� 'J������غu���W?�0P I�I�lRcdp�D>w��2�i�v���ɏ^z�u�E�rLώ]��䘺�r޹g]v�e��,�t�������_�?w��I>i�gx����ׯ�u�a5�K��z=,Ja�@LHڄ8^"³��;�\H�ސ��c�&	8�$�+0�U�}��-Yz�j��������~�2����?&�g@?��6�^|o����27~�3�<ޜ�������ʢ�x�������4��*�����S%2�ʂ�*>�U$4-��� `T���&��S�K���2�C�rX�-@.9�8�kح���pl�7�0�/0d$/�("�EBO������M��;�4
��MB��}fY\�v�뻤&!b��`gX�0���*Y��E�g\�:�>^��h�0xCX�xL�BY��.�+$!7xg��c�@�qNy6h��Ǻ�b:VE��c�zc���s�F�$�E+�,��+���k�Ν�`�����Y��ϝ7�>��ϊ�p㯽��("��'<4:2:��~*<T�����Ec�M��2wΒr�`����۶u���}��e��ZpD)1'42� RI`��j��/�^�J�W��]ZM]2C�	(�3m̀s	��E1M�`�F�����57u̝����v0xtr�\�U������s�Bn$�w���w���˓�����-ۺ/_�Rٝ;w���Tʬ�@�Yr^H�X�X*���閃�>Ë<-�M�b��%�l#m��={��+��T(�,1N�R{{}:�(�	|�@�'�(���u�B:��wX����92��=�'���C��rl��� ���fC��1���4�w�&�3�M��7oii�;���w�ν٬6mڴ������8�jzR������y�k�%��%�2��=/ۚ�lo�u �*K*GZ`cq1�ٶ�+��) ��C����r����z�,bo+PI8����/�Ku;D�-
�^���g��NI'��LJ��'Ӓ��n����tX(L$�j[{gK[��Rw�1t��ИF��J��6o�RAQ�	� BXQp����Ԡ�i�"�Ʊ׶��aɲEW_��Ι]������v�OX���e�Ǳ� '��ǟ�x��,���~��v�\��ťKOX��t&�
���X}��?<����Pd��A�i��������8N�f؊Ke	1�ż+#�38A��p,�8D��iG�U���L+�:$���؝����tHk6���
�T�1�q��W��j�~� �l~��[~�����8a9 �,8^)pឭX,ֽ����?��Գ���e���g�#7>���g���M+v�ۢ,D1Ѩ���1V;�+<�00~�ɫ���g����;z��=����K��� �c#�uu��>��C�\���.�V*�8�cz��%E�_hޒ���OZ�Z�9��d��G��[�熿���s�W��_H�x�q��x*��_ݰ��Uw���n�#�7.�������'��i�r�,���o������t��l�/|(E���RD�!M�~M��"D���
���Ɠ�Ǜ��m��s��8���=��L�٧?F5`C��|�$���p]���3\?T5E�����I���]�s2,���0�S[�B�4��|ϛ(�㜸xѢ/���M������ђI˪�k�N'�v�1v�L�E�
��'��*�F_lyDt׉��o) ���Al������e>���/���T�ʀO����������'�{���*ш��R��~���HB8�6��8f\Tlۺ���|�5A�9��e��;���}X"�2+V.���|b֜�L 3?66�o���?��E�?�W?ᔓ`����4`J/���
���x�8�Aj �X,�e�4B�D�; ^�ڭ��4U��4=�V���!2ְG2���D��J�F��F�+�����~��+�ny嵭�uɘ)r�Bxz}Z)���&�8 �NQw�,[:댵��\q�O�r��V?����ǸXR�x��]{���9"��p
]Y�29O��u15V�41S�mj�Mkhhh��lfAD�Ĩ/cj))-]��j���J�1K�CBH$~Zg��EF�F�lߦ)bg{�����΍���S`��\�� I*��������ႁ
�L�\�\��hg W�q�l�)9./ɘs��I�p�,�j<�ɦ3�����:�������B3p�/���k�lju��������</���GC*s���^��$��W��DH��y0oL5�Ns�q#Z�V��V�:�e��oh��ֽ��=�wp ׽@�\#��m488 ֺ���6��2 z����gtuե�p���⋻��gv�زe���{�����c�XA���L�ۏp7W�o~5��~%JGHD�`"Jm �H���=c�̎�N؝k֬ii�C	��qUC<��?����޹�{��Oϛ7�w��eˮ��w�n��î"⡈*pVib���ނ��1A�w玗_~�\�/ɜ�������ig�==�-r����3����~RӦ+�y���E�_m-ͺU���ڳ���w�ِM��=T�ȓ�������8A("�v ���>M5d�O?��3�X=oNWώ��J]]]p�۷o�3c� uݽ��Z�[Z�z{v��ذ��^�&����С�bؠ
3�Mqܟ�G�p��_�P�QT��!�l�����F�'F���%���������6�����yꏏ=��/o��P(!D"2%���_��#�2� AU�����((�f�kk���K"���\B��eךg���W�	N���ޝ/��GW�%K���)]��bp<�cE1րt�3d@툨�D_ ��B@~.�����=}�9�v͉y>���11n��������'>r�E�l�)ٰnk.8��w�x��-;&�@�3g����'2Y�(\Y*5<Z B!a��H-����[3�;8`��]���\��D:֘��q�5Ü���<1n`�tX�4>�G�nt�pX��XkDi9��&�Ӏ�,9��&-Z��Ƈ�ui˱{�]��;(Q�p;�0pM�/���ݴiӆ^X�hn,^tڜY������kc#9�Pw�	l*J�b���Պ)c�xs���O�Y ��Ŷn�.䊒�Ө���е��X�a�〶��񁲞�mö�d��u%�bp7,�p�e��І.:�!2�x\��i�����-���Ã͙=<I*U7>:�H�K�,��ق�������KN:�L������{���~�[�}ݪ"�~P*x!�W��V�zÒ���s(Wì��#0dY"b&�Y�|Y@�D6����68� yQ}��ߨ�]��p�衐 �O�MJ�:u�8#���̟��W��=�sQ�u@�:��ϭ���"�ɍ͞=��w�U��IV��l���}�w��=� G	M��@.#��	��4kF��ٱL L+H5rKǒ�m� �E.���<&�1�\�5kO>eͩ�l;��1Lbd�p��X��C���L��'��< �R�r���z\��	�a5G�H��V紖D:���ɺ����_��n��W�E�x�J81�k�ށ�q��~����Ȗ͛�:kN�t6�l�2@�vΦ���:� �� @C%U]	]U�O��b�
1�ye��7>o;&��fN?��3*����:;2�l�Tz���֯_�����L���D~' �pP�)��y�ܶ�m---�i�ݻG����l�8������	��'���y��{��r���]EK�5��2��=@ �}l�5G��U�BG$3�fw^{��͝�3����ڦ���R�e�/�y篟~v���x8��pj�a4�+�;��y��x�J�4lcC�,���ר	mpdPP{{k}}#'Ƚ}��c�l���	���>�����у��W3F*� }i ���ϲP@�W�aE���\�&��c�!$��Xc��m�M�ښ; ��5gfcK+V'%���x��0`M�ґH� ������ؽk�v����&tEW"r<����Q�^lb���wJ�����(�GYPCC�}�+W���^�Q�i�C��=��w�B/��
�`�b�j��dp�@�Ao����D,��g�ݽch8�����L�S	FU%����ݽ��������Vx�%-�!�;�|1�ON�Wn��@�
������8�?��/U��Jp�¢E��ꛌra��k����oln����ܱppS����쭺�zV�l���?<{x�$5�����a� 8���^���ƴYҷl~������I�)�U4��\�]\|2�tt���K��=���U�j8�Z���Xj��9������z��u�����W�c��׊E;��]�%��AU�5tEe3p������s����h��)���,��㸧�z�?{���8D�"�Y'w����g�����:�zȳD�"�zG�}AE��z[g�֜���_�bKk�xn��vtv�k�D.x��c�� 3���G���T.x��9�6~�ǿz��D�o�$]ٴ����7�ʌA��`ր���)C�5MT55pLl�����]t�{n���V5�k���o���'_/)@�m����$Ce�lēq�O�ʕ��NȐ��F�J&5�X���\~tkw��r1�>7:��W}�]�������R���Z8N�>Q�I��>���Q��?�5P%�+�n;�Fؕ�M�dA��T�ALU�1xC�*5�5nDPI��΂�jCTY�n�HdYX�l��',��']��7)i 黀���A�̡G��P��{"��J�ĳ����H�2��7n���{0��)����c.�w�2/{.k6Љ��]{�z�cʥb2������0����m�������#LM��[V>�fϝ+j)oi��I���V��}�a�Q���� Ȇiي,�~��9���	DI�oh��d�0�,Jpu�|�:�hP�.đe���T2�q}ϵd!��_�h�������XµM�W�����c���1X��aK^Tv��������+�`Y%0�,��B ������dt)iV ��ͭ�m{Ƕl�҇5Ì�А>��e`!I�TI�2�l���SO>�#=*-�����Y��V�(�*���ّ�$���кG������J%C�b�gغ�cK��� \��;��1 �Ϭ�������	���t����g>5������
�F��j����A�i�/<1A$}e`�}�"(��q��JVb��$⣅��4�L��@X��k��+���3��Q,���6o����o��g��a�a��c����5,����D�"7< 69]�480~ǯ��۵ME�-��u8۹��LS@�;��o����i��
��Ww������_��A��S릁�DZu�J�MBj��r}��������(��������+۶�E朳����_�{p��N���ꀸ�Q��׿��o~���~�4�>����3P(�ڧ���s�W]�u��`L�9��
M��'3u���}�������%[xA�6�eU�d	 �e�Ǌ����24�B���&Ο?�Kޕ�e��,x/�r�XNDmq�wN8�E�����?��w�ߓU����:j��9ʅ"�����QD��0��A�W]q��K�t�!HJ2�T֭��8{82����]*�{���(�v����C8�i���8pP���P"�&C��E�@YX4ϑ].�l��-�s�t-X6kΌ�g�mij�d2r,n����8/ɅB	��rxs,��p8�{FA�K%�w�/[��"�\nbW_�׶m�޽e��=;G��P/�eHǚol�-�v]7��tܟ�4v	��tɡ ;<$�G�<,�\V��x�?�������/nkk��Q����\n���gdd��:%-�jko�g�L�y���5�*2��Ei���֣A�uԵ���%�1٭�^���;�sZ&���uf[۴�3�y�����B�W�8�z��T/
RaЊw+(
m$�~�
�|�,�Y�c��1_�K��F�P��8� ����4��XSs�����]��X1ՠ�J"o���T2�� "�{v=��3[�lloo���w����T��q����8�y�����yh����O�Cg$?@��q�{�`p�'���ӧ�I��J����x�?�����oۀ,��m�p����s|��3N[s��� �(T+����	  0'�5��d8���&�H�A������wuu�Jx�*��a�Q��8���x�2���񘌉k%�l��S׬b����Wv��j��V(`������wT��1\T�$ �_@�{�2)t�QT���M�KX�2�Y�Ф�+φ{����:�,�j�%�NYNYadN�w�WPD�:kiЈau�;.7v^w��c��� `by��}Bб�LU���D��
5��\�wdIs��_������	rRPr�c�|vBM������)����穧F}N�m�&��ʅr\S���)�~��᳌@
��kR*�ߠƩ>Q�,�P�DcKs�TZ���9�����m�س�7w�a���}�������Z���RnG"&\�������_?ճ�%$.���1�v��H(�T6W����G�P��6t�b9~ևs"H�cK�֫T.�"Q�dD�Gx����W�I`c�TrK�P.�g҉����_p��<|�G>�W����G��|n�Z� S3*�����˃��c��n%�ɑ�B~�QUU�	)(z%�z�"��ڸ�{z^��<
+�
y�Ȟq�m4-(b(�bT�\[�~@����ְ�	KQ���+y�c���啘
�A��6���M,cd���`q�S	���ˊ"�wi��k�4Y¾_�O(	��������7������v�U��������-齇^B�;#�4��;���3�#��(P�"���z����v���ֻ�=���7󋗛S�y�����U�g���^�Z��a�\��TY��vi�q8^���୷�B�؀�� |�,��y���d��(��J�1��Q�T��=*-��'���#s�ek���7_}�}u�Oﺧ�g�2
Qi�e�}�_b)�Jyy%��1�-[~�����7Ñ@:��o�F���q�(H���xX"���z�k�'�<��i�6M>���5^MÆu.���<��~7���������CP.���
�ΓO>[Yr��	�8!mZ>�� l�?d�W�2xQ=�A�p�aöH�PF���U�ײ�M���Ƌ�8����!�\�e�Gө�������ӱ?72Ds�����A�" �ئE� �9p���#��L�\��\l�Ƚ��C��8aP*��]�I���3�L:EY�p4��N��:+���"�_*9�2-����f^{��;���h�R�ͱX
�@IEE*�%�;D#���2��n[��6c���nP.����n�������/�h��M�Ó�N�.)�TRQO�a������{��NIY�g?�;�J�����+�����(���,�88vTU]��|�1-;��ʪ7��(�2xz*�FU%*z[����ip��h8�
���q�s/�	�N�P�$�~h1q<��zr21,pyuT����X`��4�N�I��k��*a�����	�=�s<��m;�5D3�G����f�O?�����0;��;}��p2�,��,�~���@@�a����G㱪�*���R�����rp�ky��������VUQ�O��|�)�����1�������0�i��Q�"E��{�2 ���f�����.B�ABJ�%�0������gk�#��v���Kk�jՐ
�<�8U���H�@w��Ԇ���k���_�p!|
�<P�722���ഴ�TTT��������`08s���s����6l߾�+�`!@?�J�^H)X�d��M���Vr���%� *�fp�C^��>�<��=H7����Aэ7���o|c���`B��C����=�4���┲�2�%�,&̒����3Sa�;���ҹ��Y�q�v6WX]���a�#C����l&
�LkX�lymsݚ��۾�-�ɱҐ���.�ڝc���g�Yd�{��x �>R<�x��g;�xN�����cc��"BĮ�v?��X��� <@ÿ:ZZ>:�@�lappP#��vL��l^�������f�,�g��H��%G���c#�����3��dI,+-=t�`4\5�eZUE��P׾�-ǭolp�����k��D���+?n��sc���o���MM�X|������k���|0��MӀ�0c�캚ꚪ�����3W^1{�\��{�K$t�p���Q�ɦ&&e\�d�1YKzYi�#��*�ָ�88��+��_�t���E�-��cz���q����u�[Z��[*l���&<G�iZ!�&q��ql@�L�g���;s��k�{�@�XD��V�o�������{��������_�)�N��E��%�/RY3�?��O~��r�	p��q ���ra�C<&�4�y�]�\�t����z�����/�"4�8������k�mintt{�ѿl۲M�e�1����K/+jx�UW�yک��)����m��׾�ɥ�\�҆�o_q�*p}}�D	�����c"1�gj��9��K�%��UA�,b�C��z���e������y�W,==�VT��D"%�d�t����dSZ�f�g����h��Ȗ�q�[�S�0��0������Z�4�����e�`��mٺv��K.����vww�4q�=��MN<�6>
B3���ϛ7<.���m[6�b�ݒ�L�gy�DB +�t ���b#������9N�ȡCG���"Ç���za!�]�юc���vi&��,�����?$x�e�Ѱ��R�h8&/*������}��t<�����s(O�e������χNO�|��N�Ǣ%Z����P�L�R��/~��O�;�O�-|�{�+���|����5�FN� ��B6�F�-?댳.^��?�я�����&L�S"�Hh[�A�/���Y114����
˙����dHSbxj�«����h+3��9@><��S�F�w���֖i�s�M���7l�\^Q)I�X|>L�˰ߟ�������3��g�cE0&������/��l��˖.\�P��R�J��DB;|x�/�~��;���p���S$��|b!�A@nBT�O���+�P�� ���8��2�h�$TO	�#��� B�Ѵ����Js��ch��+//o��S�������rs��eX�8�6[�6�R0uNTs<Z?�O|�ߺ�������;)�A"R��z��y��L��\,�9s�gn���V6�O�� ���JI-Y�>�� rZ��L�/t���"�Hꗿ�I�}�ѝ;w�<j0�?	�"��~�^a���8C��M�J(���)����w��]R	EK�TUFzi]�h�c�ށ~�a�F����%�\�`�AQD��E.
d�46�YH�R���PQ0��x�@�x?�{�Ф��O�G���p��+p8��b7i'�R�T�����_��׶��	����n����#����SF�+ � ɲ�:sj˝w�y�Y���TmK���*]�n�k22�KF#eK�{�/����e�
�M:�^�n���� Ѕ'��>W56�����C&��Ajl��v[��\uU��sN[�bٌ�3���ys���� ��Mkml�G��rcK�O?_\��.�A�FK �4,'W����d�U�D66 ,��P0p`�s�:����??p�0��8
<V���2[�\"���Mf�;�t�?�W��8q���o��_}:8~�4��sڴi����n��fXD�Kg�\� �����h > �������;(d�H��a(GT���-!T竑$����)h�\��$njl<��pO���@l4��I�k��UUZ�d� sX�����Đicߺ@�ʐ����]��]��(��U�"תg�yظe��Ꚛ�֯[�qx8F7�m%��=���9l0�3�1dN�x��g���Q�P�)��8}{�ڎ��(�-a=�g�I��jʒbF�����pj�^��ó�>���1�Զ9������4��Dnd4��l�����=�
Z�V���v_�%��0v��s�~��_�3g���pP{��??�X۾���@�U��9�6����� �Jk.���O�|CC}���n���`Li��!� �r>�����p4�b��d���$%SX@q
�4a�{�X�i�6/J�@� �|�=rǪU|x�xg����Ͻ����sf.]����)�Mn�ރ�E�E�"��RR>崋�,�]�5��e��g.��^�<jK��5"y���=��_.����S(Ϭ����W������8�q�l����\�B$�MYP��[x��?����n2����s�nt���b�#=%�I&F��r��;�oߣ=���B�`,c��N�����o�l�|Ūko����%Q]�|�W�r�Ɲ_|��7��_��X;<����G���#j�K\���yjzS��RÃc%%��`3�5�aj ��/D��==]p���NMg�t\|�鍍u M�_yN��Ȳ��e'w=���<mmm���[�pa>�ڽs��eD9@�C�,[��e�U*Ϥ3�����;�捷�_y�e� ��L�Z����[��qy6�ɾ����.��6U�R@�x��|�X��M;�2��u5���R2�D��T&���$��e���/(B�6��� ��r0_�ZvA���7��>�UW^z����W��`�z����m�O�B2v=��}�8�g_��� a�Gh��	��x�D�ף ��p��~��<��D  ��]d��篬�o*d]E-���� hP�f
���M����?QEI7t �6r�����<�A�|�Fxw�㕦qr�'��{�uv-Á�^��Kc�#�]����1
���sy�]?�IeU,�"�.:�s֭ߜ�d fBeΟ�� �+,�"/I�)�2����¡����o���>uSY��)N�I5�q�������?���	���0��l�Tzb?L�C�/J�D��/`�A�x�ybT��n> �I�#���<ӣ-Yr�%���s�HX�(/��\𜹳.���P$k�p��%%婱8 II䯾��k��'�=��a�̙3;;;��	���]���������QD۝PFG��PPPq���jX�FJ��s`�k��}�0��X~��fx� ���g�\��B!w�E]s�u�pX���o��۽��&B$���7��T�_�I�_��BA8��h:��ѱi��[osʫJ�b^V��Xb���"K���c���}��4Ͳ���1E�bc}���p��~�kF-�:|SE�*��L�t0���"eq����,����IN߇�3l����)�%�c�B�0�N
��`�r�/�຦����  o�����'���/����G�a=ň²Hg1�#����*?�3�[��v�"��<S�{�TN�˄��,!p���jy������0���>�vWii)\U6�M&����/lM(�QL�嘔ǌ����.�s�yg�[07	'��uk֯~}-˅�`�pp��e��y�ܹ�keY(�=H�����\S����@p��ݰ,{��������N�Y�Y3��w�} �~�߬]��
��R6�B���n�Q���m(��������O��p&a��_v�e_�җ�9��y��9ҁ�>�V�������J.R��k�C��n
�����N���MPحF���ٴ��,�F|��n \Q[�<wΌ�
�i��n۾��>>ZRR;�vƼ3f�ڶyK��}�L�`H�tMg�����	�-�5�8=�<�-�z�|
���K� 9����l�x�?��	�Om����� ��!����SbGG�Y�&��g���9U���w�0[��?Q���|y$PBf!p)�d!�'��������֍����W�W�#mp�H���}��Y�O��%%�ã�8#��y���pwO���WO��忏�n�9a��%�;���k��}��=�CX؃H��sڳM�D�}�JĆ����#��򫮾��)�o!0aD��H�� ��3ٍ��I�cj���f����X�T�X�(��[���c��'̀�BV���N<cQ�&b�lב����o����X�B
{�E(��΃ ��޼��U�_w�̦��y��|�׶�{���N.��I`gR�36����|�����/�����e�w��͏?���wF�,�ʵQ����h�˱����+��B�hﾻ�_ݟ�k�*1E3'R;�\1.�l6�QL:{饗fΜ>�T��xVC�^_�EZ*�(�غ��,A��_�s��2CO�q�9w���T��4��g�����X��� D�T�$Q7\w���c���pyE��ɇ �Nă�ɤ �T��:t(��566j9������)V�b\X("��z΄,��H�O�����[�
E���t��Ӈ��tw�`"��!Ny����"'X�x����̙+N���+�Qx2�ۍq܇�$ocK<�<�?7}��y����˭��|��/?�d"9JS�c糹�T�@�g�Q7��jꦜ�b1�&�:�v6l�444����$II����&ŻG�i0�,h�z�Y��Lg3�L2C��]�_���V��ϻ�r�P,��t��־c������ٱT�g0�ҭX����"�e>O����A���0��"y���!�tᦀ ���S��x뭷���g�4'<��G��У[�����ND!��<�̳���._���/�1�}���]�?����TI���Þd�k�>%����s��g�iB�⫲!A�a`�RG�Y�ȅ��2�,)����VGj�ޗ�z�O�SUUi@Qa*���
!/Dcp[Ul���8�~P�)lT�M�k��(윹So���;��~�i�i��'mM'��ٳ���
�"2K��\2�RX9��Ύ�4%B��\���d���ݎ?I�OX�Y�q��G%Z��_�4��aEÂ5�9����3_}q��m���_4����0�Q+�͙��R��3��3��aUII�����Gx����E'bS��xp��e'$���!�i�R�x�QU
 �]����{����ۿ/$��ՕB  ��{�9�������s�=���Mn����5]{� �:::�1�|)�1{���?Л˕ζ�����������|�_���)3�M������^6/
��lc0�u�0�x �(��Fzۖ��]���VPD��M�����f�_])���kN�'� ��&5ߎ�L�vӱ>��G��Z��x��Îi�8�"*�:`x�������y��N��i�/*�_�ж�B����
L���`����2'�G~#H�p.��P$∪*�����������P�1^�g���Ka_!;���1ǿ$QbLcܿq'G�����<�sά���������$J#���=唥��
���$�e�YZ"̜�`訩�*.[���j�C>B�����s�\OO���H"��DµՕ�kV1��7\�忽�w�<�̡�HPV:�!Z���R,��c?�ɎX��P�S�����(~v����ЕW^���~w�ҥ�� {`!6oޜL�!���GuIi�M~�����`>U%��pD�_�xT& �&����SCmz�S�6��@׺����Ön�wp���]=��}9�
�(U���8;��t�8�mkRE{~5`R��=^d���z&�iN j\�f�Cyw�?k���׭�>}zwOǻ���͛�Ue��c���ҩ����D**ex��B$PYY��)_ 1�C��W��Ђӡ���50���2��������S�C}�5�7��M�q�9xX<Ӡ'X�r���Y��2����EY��
���	�K��c,۫���9�7��۷��g@U¶�Ae	�r�Ej=_����4g�֭o��VC㪰J�8���dGʰ�8ϵO�/n���eQӌq�)^W'Į|�o`�%��X@l��[��*�n�41��7�1�����S04����Bx�Ϻ$v�q4�qnB��scF�>Ҷ��ݝ"x���,/�1s^}cM۾��)���"�-�����~d,���7���K��<�B��s�pi!���d�O	�6"�v�\|J���M��t�����'�7���~��GT�L"�O �J��G�����l����u�����S�$�� c�H*6�����w���P��0����6�Qd)���05�����C����9}�W����3[��5�`�]�A��	��X ���ֹ�Ɖ�g�c
r���7�>�g��/ɮ�lm�0,'��َVQJ������p�="�'b�w�H	�V&�U'�z��鴪��;?��e���yIQ!N�S}��PN�Ӡd��́($>��9���׿}�������x�i�T���̧��p4���XB/pђ2l�.)�#�B��u�~�߀��9��(�&i���aN��h���e-��[S[v�5g��Ǯ��.ͦ���C5M�8pH��n^
���v>��;.��L�H/�; e2g��������'8w�[�!
;10F���a��Hk~L�C0Y�p��S?��[K*�<m����m���_<�L�m:��h	��������t#��M��:<4����r�����˻������l��5�AC�%�3x|�7���q�{V�~-V�rq�¡X��fjn��l�Q-�q���h�[�T�a��r�y�Ŋx����b��1��~ 	\��8DXQ]u�������N"M#Êe�Y��I�u퍫V]��GS��A�as6�Nea����?�УO?�L&_ 4�Nq�͏O&&�Q�]+�q�#lƾ&�o�#����ev�9�e۞�Ͽ����+���_������c�B����a�Q�������Nk��C�"]�������I$5������
�^p3�B VA�r��r��X��7^߷<G����~=�b��iY��%S�c�A���?��ϗ^vEUU�t��O�:$7�Ce6��a�Co���(G�Y����s��}�m�C��!������>�{"�s�ke�[y�X����O��;�ih�׶w�w�0��'i_׿�"�\W�L���p����Ȍ�W��ʷ�8c�`�t�����ka6��x��I� �V�C��P$��k�*��z�Ȥ���R��%c~���'�� M�*�͂��r}C��΃x�bD�G��#G�jjli��@��p����Ç;;�)}d(�ol��غ�(�0|�<��l6;��S�Pwd\]�qBAa���Sjꛛ]�_�f�3Ͻ���/��g�=eي�s��4\�������E�P��S��'�^EI��F<ƱBS�Ԏ#����bQ�������F��W�\��������s�=����bqXI�r�`�<�~l��ı�?+B�kZ����7�`���p�7�u�]uuu��`�Հ?޵k��3f����F�#3��&@�U_�X]]�q|(Q�¶`YG]��F�	r۰$#�2+qX �1lY���;�A%��:E�ܺڪ9s��;tpGۮ������QIl�R�`�������7���=nQe���cy������7�!�w�t��u#����]p�y���!��|������K"����s�+�|���;vQ����S:��� �V*K�3��c4�-�򊓲�B�c�j+�4yN�rK�p�!T˨�2���~>���[Q�fRUUU��ٵ��m[�Bfdx �͆#��@�4:B���DK��A���m �t-�O���ǡ&��!YQ�EO��kY�D,ֶ�-�%%��6�$2L��9۳'���)G
��_�8��\�U Q5\�f�.C����
���>�X<�5��ˁ�a9 �ǁ5�����6�ଡL����S�YiS���x����Hƍ\NfUn���
�|��}�5���Ll0�)o��� /W�{�y�	��8�
�k.��}���#m[^@	�=o�6�ܞ�~�㟭~�5pa~%ʭ�I�5���^:1�(ؖ�r-H/��w�t�a:�ڏ]�s��'�������-`y[�8C��r>���$|�_�*�-Ь��^�*�ՑAL���X@��l���(PHJ�[S�"J�p�����״-��<�'�*�6���lk0��֚X��E8�σ�m?ҾnӖ��<"XA(���kf��d�F�|!�d�� ��uz3D���s�z���'�j{{�;�S�Z>�,+�a����A�|������i�,j�E5z�E{6I�͖��g�iL�2d�x�y�zG�ӟ�[���{^�2,��W�SℓG]d���R����/� �������mK����T2�	���2uS��Mm��/Ă^-˳hV����cό�&$�F��d�>�f��[��(棉���3�Z����'������*j����d9��i|H��G,�î����������+��
�EumMEU���e����(֦�v����r��sǤ�� É�cZ�k�5�iq\��y2��N�Q��cIМ;cڪK.8}�)��(G�P<�=���=�"�c!r@��r���\z�TC1���f@m���TTV_xᅦ��(�H+!ޣL�vxFr-WTprأ��<�w�2zZ�(����[��U�t�'��E\rw\_����������MOL���ϸ=Ξ�/���7��V/\���@0W\~��E3��/^<2/)�Qp��hotl�ȍ7\~�E�.�s��$�箮.?���C�m$�P��@�>�*fFt��r`�d��h)��V�����?㹖��c��ރ�FɆ�R �==�ccc��KU�$�3���q�������`�o1�M��V�T:�'����=�؟_z�YE�� ͽ�<��+����A����H�7���<��3�:;C��C���d{ a:sT��DH�Y���\L�3�tS�j��x���7��(rT��@��mm4��	`Q�6t�g_X�~�w`M>q~�I&Y6�ˍ_�x'�C�B���m��4m��`mL���s�P���*R�6�|�0�f��r)�s�䲋5g�tp�`C�5X�Ga�A�hp�"�͝5cZ�Y�6�̽�~4��<ᢋ����,_��rp��1mXQ�)�W�Uz�NEw���k��2�]��px�e---G�v�<���h��74�{��WO?��k��q���<�������^�K(X6
ߑ`R�O��Ȩ�@�'`y�E0=�	��M$���.C��
أ>�����7m��{����S�E@��vp��657B�J�	����_^<�
���s��)`X�;l֙��8�M�z>%Ë�,Z�`������Y,+����YS]u晧�Cݰaa�e�#=�#X,�
nx��ST2� ������K�eӦM�x���-Y���uziYe$.-�6�5j�N$}����:8�y�tJ'�������1�Ij�<A�`� ޅo���(EF�c�� �ZZ�̙�5�ٳg�q��#��EKB��y�_	v)@|iA�"IH���C�ۇ�u��������Uԃ���\A#`XPH���!c��#zs:Mk��_�����9	��$�!3�Kf���}r[�h��,�`��p@�(/3���`�B&ܳ�u5睻��SO���$�Ά���7�{��^jo+�Pl�����ǵ��(k�&G�����^g�Q,?���L�i�<+�?R���@!�̪ReMYY$"R���,%z��,]
� �8ӢX�]�YHņu�/Sy]����wcci��L6�z��E�>��9�l���;k�}����{��_|� Q��o�=Z�8��I�m(Vyꩧ����Vhl]��/�й�^{��< #�L>�[7�����?<��pi�ʫW�T0晲�At�J�	ܶ�^�0�������C��z���\���{�we3�$*vq��[*��8 �|��oi������fߧ Μ,?�DS��SϽ�h��sg(2��2����vm����!�k����̡@�Ӗ%�7:4����k����`u?=|����{�7���糐�>��cX�8�ܛn�$�`;��s��x���"5-�s��d�������^|�iV%Y��V`�4�b��8�7��!��8őI}C#h�p6�s�$˼f�*��*1�`{�H�5]�J�3)�3���p�FG�e1����b��0 !��KEO<��%���C�ňY�TÂ�7׭}s߮���@�϶\z8����)d}ĦpM�8F��C�l8����"�-nf";Ký�����b�\��u��c��9�����X�G��n�k������ֆ�(1`q�2V]�%\8s�Jw��y�����y���ll�����;�#|����Lnw�2�D�*�tӶ�[=��M�3��iڅL��E^�mZ0]ʲx�� ]�aZ��I�d�|�V������f�HM��:`ŏ.ޠ�������(Zu���5��g�/���ќ�34-/�L}]KyY��*+J�vw���׿��_�&���.\��:+[�>`Xvwgׯ����^����(ܡ�����Er�zۣQ&��xp�AI	s��<O��f� ���;{�w�=T�4�稍�3������FB�@@���l���V�N��!�����t�7Ɂ�$���pq�Q��\��N]:B������Eb?�TA���n	&8;p�# ��w��$��$�>	�ji�849ğ�C&�8��s��������n�J�ӛf>���N�X�pDF6�A�4��e(��f�;�?����N0�.�"�f�%�×0&��D�{�-�(��|���x����Q�ӛ�FƆ;zz����3gΜ��=FȢl��K�� ���� ����`}���~ֿf !�rI������@�H"�f��ҥK?�Ϝ}�Y���{ؼ�"��8]��4bXF�D��f��jڇy���N��YΤӡP�*�.,Y6�"�,mmmp��Ϛ	ot�H�lA�=o�mw|f���?��x<�]���A/�y�E�O�"�F�p\ Td��>JG�"&��8��|�;�g����ذaCUU��_L�]�xb���g������g��U�3�H'���31���ї��Ű�Ř)6�i[+z"CIP�J��]�쥗��ٚg{c4%�ח͚Ӵi�6���$��"��2�(�<���c#�c�]�kP$������8�f͚͛�"�f��D�̝5{�<^`�ݰq�}{�H.�X"	1���>*��q�ڶ<�qP��#��_�����p|c�� ra�k�> �^4Z
��$R:48/Y�lYI����[�v�,/�߿�
�z:�Жi�ye�Hǈ�����g�3�-S�Nm�R��*)�NY��&Mq��z����B.S��XS^^bhIB����0�_���"�bN
��a/�:�VEi�o���U�eR�7׬��k�t�H���k���g?7�����L�v��N]4��$���8�5ʈ���]���x��E�cP6�yY4�}
���}8¤/��Q�P"=��֘F�(�߱��l:�l ��H�*u�r�}L��I�L���c���կ�^��/	@�������ax�2/ntww~��_)�޾U����'`��`.*{'���2"(�� �hVH��=�؊%�O9u�V���z֏Τ��~w7\&bE�E���(J�w������}�𣯕�DE�Ռܮ����C��d}����d����c��%����˻C!�ّ��=�ܿ���#�X�l6��.����� /ɕ5��T���?��O,�2H.lh�e�ݼ~ϕ߬tr؞�R��wm���/}�_����]e��΄m���B1���� ��|!�*R�ȆBe=]C��o�}��G}��‐?ri��sM� �H�	��F���UoniI�t�a#�h6���F�"%�#�3�<���<��u����_�{� 2����rD#-dI� ��ӈ�O/�!�*���_Z����j�=nW��橑H�p��Lpآ���uS��,���������hI&���s=]����d,�&	ż�\z:L��瘬�^�p��` �+���2u�体�pz&��ӝ�=/��j]K��Fu��9߰aV���8�I�͒UY���tl������p���u?���E����{��, d�SjB+�8�iJ���h_O_댖�����kꫯ\uQY�
�d����SO��6JDﾵ������O�HT(��
���.Z�S�Ř�8�.��1@������z𡎁�����,�,��?�3:o�9;\^zdߞ��J�"��d��CeX(}If���ݴy3�i�<p���N�,|�m*����X?L����, �k�gS�^{m��X�W��o�I�	>�>+E�����G~��_�����	��3l�u�m�v��_������^�"Bm zI;�{�lSi�رC�xpq�p	�\�t4���ga�.qk0|�Pדyv����h�@O�`_o@�E����P ��ڃ�W��>;\�-혲X���C��N�^E4|�i�O=my�,P"�-?�h���k6m����&������H,;�*�'RqT)�`�49��P��A�U?8���}O{�q�3��%U��i?�#5b�(�-��9@0�N������<r�������,�u �_v���ڻw�aX�lN���;��z|ߒˀ���
w 	�2� ����K�`N���t"nh9���`g`�]6���ع{��}`,���h���S$fޟ� �Xd�B�����+d'���	�����p!z�6�h�(H�G��Ga�[��]���W\q`0% �1���C|/������4�!�d��+�N�B?�
�aW��Hf�(o���S�Z���{�g���J`֜�-S[UY���{����5���.�77�����ぐOGMp�q"e�,�x�<e��.��6FN>���g��ӻ~�h�b-_�UI+�l��b֬YW\~��|92߳g��� ��ŋ�VTT������?�,�A�y謹N27p9A�1U!Y��hZ~dthth0XY��#�]{9Z���z� s��/��y}�"W���e�%�F1̪�` O����&D��K&}a)<؛F����_�c�a�Fd�k߅]QY�62�3:ܛI�uw�j.�ݲu;Vo��+��-ۆ�3��h6!P�H���ќ
��Db�;o!�?�C<�r>� �L)چKT����f��3�.Y�������^Z�z�HlV�@b>��TV��^^Q��;v�-\4��1N��s�F&P8�112޽��粹�K,nh��7�e����D�[}M����NX �-]���sχ��]~dx�����ef���HP��I'��A4��"�-`"��/ߺ��O���\v����E��;s�������FBc$��\�1<�-����d�]��l�d\H��d�AK�.bU�s��(L�塁�J!n���g��)	�$�I�B[�z�����ydr��8� 1�|"��r��r9 ���ؘ���B�/�Hp?^�%��X���uq~�� k[9]d(����n���{ĥM^�h׀��'��py+�,���Xp�(�Q����;�/r�0�`O��H����u�ֻ~r����̩�,�<�Pgr8�x�M
	o��,��(����Sױ�|çfMoI���x7]˓4�����5�A�2Ep���"=�cJ
F0Z�x��gE��η�u���?��ѧ�|,�NHrAO Y$;��j���'�҅?�15oN�g��q��TZ�a7?�@[�&ĵ��4���-�
�t���˟��tKKK}u�(�Y�J$�P4���}�0��R?ph��s�/�}�y�Ƒx��D�u)Ub�����ie�(S�h^Ie�:o߾����1m��P���k:|�pA�,Z4��4�m��ѡ�Yg��sϞ�`�ۏ�ٸ��,��q�M��,Ǔ�ȣ|a^Bb���|�k_�?A"�jo�l��<m�����D,Y�e�P{�0�MM��H,6�uu�)�]��/ "l�2���ea��O��%���~��ʒ�+��T�
�I\�}ϕ�����ȟ��~q�����m��C�'6��c$�*��Mt��x�[���|�M�M��>��`��zt*�Z�؞w�%�~��ߋ��8�֊�����T:QRR�7ˉ�_A�k�,r.�R*�|���}�Ϭ w
0C�u,�$f]SGưD"�"�D�2B�M��=z,�����L�'���'����0gޒ3���w���g���7nnnn�����L&�1hi��t>��o��Ên��0���q����f�N�|�!w��P���X�~]������?��/_�Ld�x!V�v���_�����dS��b,���X�v�9;-\��3/��w��^���\rI��	}#�1�g���晐'ȍ�w�db�����
����c7t�F�g��{�O����/�De����̂�A�C�l������i5������ckA~�w�0���x����G���ɥR�`֫|��y�O��8x� �i������/������l2ô!n�s3���H���L�H���8�"�]+���Ng9	�y�5- ~� 8��5Z���󗧟��s�LMuy�������~湥K��[�ri	s��(�䁥b����d�o�tR�P]���.��,Q0��t4�������Z]s:w�w���#�L� ��;�lܸ��w׫*�h�lS�ܲ賽�����+
�P=l""���H��=���`(⒉�<�I����dɲ[���SO=���#/�O�2ar�da�h���Q����Xl��]�CHJ��_�p�_��	����	�_�k�74��G��[�Z$˟�5�׹����;�\�s�wߚ�+�
���#㚪�7�OH~K�57���r��ܔ)S,K��:N{{���>
��K.��{zz�x�0�����yē��=1�'�(�B�J(Z+��Dˢ����m{�c�M�beկ����կ��~�oh�$R�w�<xz��HXo�f&zm�"+�1џ�c���r0+��ԧ �:���7F �����B�%�\y�֭ۓ����ep<]VY�7KDT���
�Bچ��(�j:�I�ҫ�Mq��-�$u �.	��U�����m۶L&��a'���~�Кo������ٳ��f������|�0x�u~;u��Tgg���@=S**�9��+P��� �|]33C��p�ħ
o��&l�������w k��>ҝGfF�o�'��Ubl����n����Ah��Z^{������fX��3�i�o p�(B������aJcSCs}m�ZV3�ƛ����~�s� -H��ԉ���x�^T�6-T@+/9��GE<fK�
����6
���8�
H6Ե\|��ʊ�G��)}����R�I-������6��fLmX�`V&�~��
���a-�-���٤������sg�n:x��˯���KHb�P>����+ޠ��R��8e�����_x��D"�ͯCVĻ~���~8��1����Y��9����N��ǿJ��_�����۵}�v w��0�����.�����[e0�YZV�%��ē��Z[[�}� ���t��,Q�Y�$�Ă�T��@�7��SO]�s������$�c��2֤\?s��[��B@�<�g�������fLomhjjj۳�4�����#qǴ�y�����;�J�#A�F���j��B�P�(����jk���6Ü�
��'!��$�DÑt&���. ?��i�l��#���A� GSO<���Q%̂�e��D*A&	��!8��D��!��!L	��{�0�؉Ϳ��5�
G���n-�	�E�[)����W8�� 3 �SąҜ������'+�J2�uH�H��w$՛��򢓂7�\l���K�
�)���&�j.��Y.6������-{`EM��s��J]��B��yT@$�O�~�a�4"s�G�|F5�UZ�'n��e�����'���7L���z�T�W���s��g��\'8n���]m���i�`(�@d��d& �J���۬���j`�P6�u�&<�:q|¢=@_aE��{ۻzk��'�Z�p��>x.�˭[7��Dr76\;�/���Qi�����)�@���Yrlҹ�QU��4+�1L>��D� \�������WT�����G��c�[�Q�&�IVD^ݴ~�]���+V���+6n(-)��b���p9��� J@��%h�0�~�Q ��������GY�s����7<��������#e���o��ֻ���1W��윤0�wΕW]Fx�, �p����}��m���z���\ο���w�m��B$_Щ`�?U�il*���Gʃ��q�TCk5\���sfΘ�����o���O�rp�%YB�����:�I�;���R��.66p9X���L.;rŢ�S��Y��;����.��ںj�IC�����o���Ǎ��G�G+��"���3�]��G� ��f��W%�0 'F�w���3y��g_����8e	�j8�L���b���A��'�Ċ���*vA��#�B�!�`Ǳ��hߛU�7C�����몫a�^w�uSfO"Ɖ�S�P����'>���dBD��_C_��/?¾�K&�0v
��I�+��������޸i#/ *�E"�3Ί����?�w"7�����Sq�@�DH��4Z�R_QQu�ퟆ[B�:��������{]s�5~#Yww��/�Fm�ԩD�������j,=��P��!#(��p$�\f��sx��aޜ�/�z��å�u����?=�؁�a.��1(R<Z\�727�|� G�_�z������f��W\q�ׁ�~�֕���Ã�:`Ӝy��J ���@,��L�8�`Ñ@����p}�p�9#����)�3��E5�	q68u��1cƌ@8q`�ޮ�@�Ӧ�h�ڜJǟz晱�F��9TybX8�;v���:[�ϲ4���`���6�%����m�ӟ.��SO�_W7���j�"{v�J���ñ` RW;%�,�#�e�Μ=���IV$x������!_��~){d���'���v�i��zǭ�-Ͱ?��������YU�hyi����4�R�>��c�=;�t,Zr�e��OWV�KR��+/y��_}��XfBs��^����c��,�f4 UT(�]wieyx�o������޾8G�`1aAt� �		�e������g�u��x�d��gV<4*�"��zoB����O׃�&�Dc�U�~�_�?���W^}��uz�*�4�A4_V�~�3��x��mJ�0�,�Y����������8%���9Tg�	��xn��>����{_q�P㒓֭[���U>�qg�h� rT��	�i�l����|�~�ѿjۓL��� 
(h�H�$�MN��q<��`�Nmy!D#���7W����F�X*W�H�u���pC ��󨱐C��ϥ{S��޾T2�n������ЍA�L{�Ĭ�GCk�_�sL��ʊ�\���q����j� �3Oٺ��qb�+�m��B��x�0!�eX �x��F����N��^���vc��S��l��r��#G��`8�I���*B!��>����g���C��PW.o�ܱwp(&�L�B���|�쏤�X�±4�����3��^��y��I'��(���*K�K��.:����d��#SZ[�?�qӶ�n�siʴ�T&g�)
lۧ ;g�������:Bz~<0�; t��K�9�iӦt�%9�� ��|�� ����Œ��UW^���<����c�f�퓝"�	N#?q[�7"F���-ho��������DW"���Fs����������%��TF��d8��7����8x� /p�䘟�Q`}	=?5h��%OT)��X�g9�u&�d0kWWSzժ˖/_�����>�r�@/��a	��c���i�Dr�/I��ٞQUQ>o�K.��op��?�>�L9��Qb9�BjX7�D2%Kb<1����ź �}�F��x[] # $�6�5o�ٲy}&�#�`OT\`3#7)�Y�K4�x�]L�L��$&������W_Wo���/�ygMUվ}�����x|lddʥ����������SV,� �,���k��CAT�?��(OPP0���g�����/��;�r����8��~<�!�Ν;!>�={v��$3�����)�ɜ}�9��wϿ�ۿ���%K��Y~*�x��h��(2 �</
9�t��"0�LA��C�G:�a�/�w媋*�*�5�,:P0�7n:xhbg�Q�c�\{|�O�¡�����@�V����r!OS�P���v��-o�ݺiÆ��;���ϩ��1�$�>wvvB ���A��n��?�p��,��`@HU��E{|Z|�['�*|�. W�(�`�\oO��s�;�c�|����)$����9�Pyx�p��#��{��I�����1}�U�j�	7�M�&�^��e$I8묳���X;�v��	�����g���k d�Ǥj;�l�%�6؉VG��o���W]_�25pp�w�=��ˀyn��������z�����/�<�C�h�6�/���W�>E䜖��aJ�'?u�-����{{��C7_u�m��������9�4Rэ�]�?���4�ϣ^�?o~�o�`744�	{衇v��5cؗiӦɲXYS�bŊ�7�T�A���{3�'?т�`jY8�Yb�h?���0!8x�,�8�ZUTU	�Z�j��>��������ΰ��j��9z���R��$�wѕ�b��ɐ���Xhr��/��G������`�$�]~�٧�vv!��s:�`��F	2[x�r�L&-!�%ԫ�����~{{�x�k0��Sn�8�;ɭ����xüsu-'��__y�������@�4�F�H�w�۶tu1]a͛���=�*\r鹕e��^Zw"Z娣*�C����()����-�6gN�*Ѯ����4-/ZV]^Vc����(3[�0��+}�����㲪�2+"q��m�PxT4�~xD03�o~�[�-�=U�<-ZR��J�6�)-S����������a���DJo�X��п��#}��9��,�A�F�!5���>����	h�̙tI���e��;9�Miy�cx8L��[��ep�� sy�q���o{&�'Y���M�)h&�M�a"*c.��DIG�  ^B�b�F!���P	��y�G�
�3�X��
ӧ�e�	����Ғ�x2Wa�e����B�)����Nqg�+��}�O�V=x�T"xJ}��+��p(k��l2�r	Ub[Z�mS��}�UU������9PE�H	*�@DڄYѶնu:M����h[m����[�6cDEA$�
@���{7���}NգD@a�_��*��{�=g����۶)�Q[��t�dUry)�%[��#���eU��N00��e�W^~�w���Ғ�=������ii�"�F�s����}�;���v�}$���G�����d���q�O�����7L!)t,5��=��g��Y҈�[. ��Ǣ3����jpI�
�+�]��d&����~�����2��	XfE��t��{44Xdp�	T}� ��-�U������ܵx�b؊^�����>�u�`�`���KK
������L0��"����̛3v�(��O�z�/ڇ=͜���)���P�C���Ji�Ÿ$��3 d0��7�����ӧM����M#y`Cw_ye�(���*�pK󫇕�J}}}}����xa���gr�!��+B:��������K�nk�9���eY��K�_�d���e�@[W7���nY7n���j ���>�z�kZ:l ��\b4��O �{���[x���O*�oik��裏�������!p������N+�hz�vXiuU���<'ñRd��H�m��7t��]-�����������f@����I:e�N��J&dm%U$���C}���-*,��yy��_=,o:������@��ʋQ�а�>�K�ӆߟ������_~�F)@�d�5���R��3j�㟞~���X���� ^"�}��������I�FN;m�~��cǏ��9����w��;w�%��N#���C;9"ԑ�ecَ�� `���b��ag�u}{�G���)��DQ�*e�EE��(��r/8)Q�n����}��
^���t�I$�56����X&oa���s'L�z�ܳ{�k#�h, ���PPu�D�y�������;::�z�)�p˴�+[j��6����OK���欨�eA�N�	�J�����.���U7�8f�x=��0�[ش���9�,��/� B�U)�$�%k�a�R�;����[H/Yr>|��s�m;DA���,�f��a�G�P6��%B6�<�'��Ǡ΂�g\u�U�y��^Y�[~��G`�����RC�ᵽ���eee]t��A� �y�
�o?ƪ���Á��%t�(,/�E�(*�1b�����{�~2r��`iŅW�8�p��})AԄ<v�%<���m�,�$��XIy7C{�)�T�����3�lڴ)���~8�@ǌ5f�8��k֬��e��ap�Ӌ��ŉ4�G�>����Gv��	���Vy��p8:�Ɩ-[�HiqqqA��� jj��<
8��@pP�ŭ�� �ƐY`���u���)�������;o֍y��G���#K�r�0�+�L�$���$K&�sMϱ�}�{����F�([9 i�wOݱ9z���h^��q�˯���Q�P:�h�q#�`� 'GM&����|�����3 �S�ПUJ�)�e+/]y�pH�<ñ5�9��**GO�Sq���ʲ�2=��2�U5��
���=��c��4wb"E���C=:|;;����P6n�`�����_M�z�<�����qGwB�|z:�V᠏o p�t�s%�S���SP���_�ĝ�z�3�T|1ۤ�Q�T�e����NM��$	��+)�c�B�^�҉L��DlC�\+'H&S�'��+�mEy�����iz� L�F�'�0-��q�`w0������O�
>s��P��Sp��̚�x�����&�7.��ĳ�i$��KJ
n����,:+��kh�����=����K�Q�9D(�!13���a���#�pR|
�@NӒ���?��w���9|������pXTP<2�������[���(�6�o��:�q��鿯Y���݇�H�|
DE��<A���f.hha&�rlw����.�d�	�퍛0��������Ț�����]�\�񹉸ʭ#w���km�}r�S�iA�B*�ف��,J8�~�4a���ͻ8�{�LF�z[D���n���p�ͫn����NIa�aj#ƕ\y�{nذ)�ѓ�`z�A��N!��n��C��\[��$ѻݿ���?f������/>�f�޽��lm9��Ҹqc��h<���X~�T���-(��,���\��DOA�*R{,;�!�dk9� ���D��wWǡO6���l[G�(s.��5Ҕ'���JNn�JY�H��d��p������F9`nv�g&�0D������t&��t�+T� �����	��v�ȫ��f��ͤ�]e���8X��\���55��#k��^S[;��իW8q�ZN�\(��d�����U�9{�ͫ��1}J$�W����<WOO�_�y�-[|r�%�Ϟ��K�WU�$���{���S�+@w��G��x)�O�����Y�x�����[n����2)��c�R*$�΅C^Iq�n��E�B0�iM37'\ܶm�K/����B��Y��
(X���X�x��NOg��������M�F���aPa�ihjܳo���עEgT���k������?v��ǒ��mZ'�2M;[�.�m�N`**
jjGmܴ%���i�M�"S���������ݽo�̙%E�����S��S���+9s���cƿ��;���ҍ"�q����ȣ�6+bHQ��?����0~�I�7|����{�7M�ɥ� V<lcc#�I E�{��9�G��,5`3Z�Jl�s���}�,��U,	 V������[o�y����*� É$W!R*�m���i��si
��>��5��r9��poO;���˖F��~�Pc�ATV�)�S6}=T��F�$B��#�K:_gE���\R�TTX
,h�ɑH��5>ݺ]�X�\sMEee&�njjZ�v-X�W��� �0�hV�����V��M2����W�X����Q����jع;�1u#�w$�#�\�5k_z�7���\����r�=�E���A�4��9p�ׯ���!	�����W��*zἮ������{�'�4��C��iCU�4'K���@b���#srr��PX������G��!؎zF��V___T��bŊd,V����YQ�
�՝;w·�u#IK?%I�5k��+TUUq�ZI��gK�XV�e4������{��MK��.\���q��1jz���l+�6��YneeE,ڿnݺW��bc��bX�ʷNz��h�%�qL�b���@��0�pLL"H��==�]�����1E���ٶ��,=��J�F�`��N�@�b7j�x1���`/���LMl��9��N�Y'$�GH������}I�%�1��~N����+��믽v���L,u�_s�}�.�6ENP$nՍ��|�*�6��l�����[:z-9{�j�Z \s�ս��c���u��|B���Ѫ�/�9F�.
`6X���6N��x!��{�W.:kAOO�Ï�n��O���*�����K����U�;��o���Ç	����q��_L&I�S%gQ � )�#��.s�cV�	<�S}�D������w�eΜY��~D�2��h�d��0��k���m�E�U�L�����?���f89N��Z�V�]��eZc�}��W�Ii՗LD�s���ڋV\�͜ɭ}���[��SZ*�߲�o~���,��jz�5��˷G�;������M�x(��Wdd�'W#lʲ �L�8�'?�ׅZ�Q��]{�� �I�ՕE?���V�\��R��34�AQ��ѓ������ϵ��4�C^"V����C6�KM+,���D@UZݦ{��O�L��ƍ_���+<Nq�(�~�ӓ�H�fd��6�Ww�����}��L�Ȥײ`����Y���rpz	�9נ�|0��lݠ!^k��_()*�馛JJKa3L�0y�ĉ�c>�  ����u4�4 s�E��%��.��ۺu��^j��e4�_:�Im[z?Y0AHjS[�D��A	+������0����/�8Iӹ���=��v���������s^(���ɖO����>�r8�<������ڃ5
؍0X�0N��@��i[�EX6�'���rr�p�ZVZQ^^�c�XP��L*-p�,��&�ڐ�>������g�@n2�=�p�3s���g>�;f�SQmS��drd��_���������5d����g��aTU���G?O�ބ�#����K/������}��ﾻ���8 �&�@i�L���C����f2�$q鴁���m7����'��w(�E����T�#��?�w�;o���?��h$��V�����f6Eem�h$PPX��t2�L�cP�Z
B�y�Om�����3u@¯~�Kx�sϘ����.��q�=|���9I_��x��\��2J�(�=q\�uW}킋���?�>����--A��z:铱Ul���3�h��g��xi���9^���L&��5vP�P���
���ѣiv+��3u�94こ2�M#q�8��7�z7�t�Xނ�6��/��NYe-�H{{���׬Y籦���u��"������ ���w����	���,q�f-�M2v�ؒ�0P�wl����.��w�3f�Xܫ��H]���cd��V�K������ʞ��p�x<�t6!<N[[���L����9.F��) ����~�����#���EĹ���D��ؾ�����y�O�X2��/���E��y�]f��G��I��N�>��::�{�= �˖-�_y�s#y@~�t��54Po�g��a���9�a��f��*[^tN[Sӛ/>_3r|��:at��I��/�����འp���M���h�Vy�Z���b��p!�yysg�9��sr�---MMӦM����-����i����t�,@x��8V�&�OX(A�3z9S��|Čj����8禃�ڸq#/1EEy��,w�������֭�~����i(4-���t�̙EEa�ӆ>u��?���e�!	Ŧ&���dLYx���~�w��L{w/p���q�X,
7��>X
β}>��qK��.+)���$��i �e]1.�I���/p�NL7EɔR07���7�i˦Y��3�n�'���l`yI���t�W
�r�	0��g�?C�}Y��,ڹ�1ra��4�iL_,	��;�z&i���(�>@���e,õ}��*9O?����?Ks�͌]XX���}��ɜ_��+[�	k�dҤI���ǎs�z����������͋F��
�.]��q=����~��'��LN~����p�W]~yI�ۈ��._���[�4�.ˡ.�Lȶ¼��ps�gy����o�v��o��&z�_y��Moǭ�s���t����ǡP.���S�yz�U�o��W��s��b�"ʮ�B�,'QRWMrT������0"�٧ϼ��;杹j�E�>���C-�Ux��0~�%+.���[���"��'��[�uG��Q��ޏ�v��ȼ�N��E3-��b����v2d�����[n���PN����?�q`�a�0	A�n�q�]w��-��2L�7j��W�Ys����;���Cݽq,C��f�Ӊ�G��bZ�\�_{��+V��3L����w?����h�_�o���+��
�@y����;��߿o�ڋ�-s7v�-�d��-[�Ɠ��dq����=�g�p����k����3�/9��wֽ���wL��F���$������Pn�m{������?XV�믑^��iS�,_�|�ڵ ��SYYY[[�	98�P(H��Y������io��o`ٓO��5�?�!��f:�M򕕣pĉ��Hz8���b=�$�	}�6my���^[��̘J0���$�(9�yR�qC+�i61�S�L2�!(ˮ��Xo��y���]&��l6*h��{���~�ȣ��̙5���8s��啘�����Y\7n�/���v `��p�N=203�I��[�ɬ�)RQ�*S��xc���#�o=�( !b�rj�C��&�.�ћ[[ �������n
�?��������+v��	#��Ϛ5?O�}!-i����LQ�b�t��/\���ػ��5�:���]K�,�xU�,E	�u�9�率[�p଑hϲ�AEJ��8���5#��ho�~��'��;p�u7���$$��5$Q!�既�|U��(�U��Y��W_���;��iQ����/�"�L�� 7۶$���u=i�i��5Z<�>���;Z� �����~�pQA��޿�����zj��ip�+V�����x ^٩������"���C�;j�+�k�y��!�s��D�"g��i3��T ��xj�ν���ېW�v���n����� �|��u�v��NZ�d�DY���A͡jr���\�3�U@�`��v���W7o�>z��^ [���>����&O3a̀-[��������ˎ&%�Wp�d�ʦE@T�$+�Na$m%��
�!�^&���d�7�q˘��2��*��~�łUa@ۖ�-��T~�>��O��z�fe��0۱cǶm�Z�ZE�;֜9��ز���.�}��?^iko�/��TK�IN��_�@UxU$�3��젇z�4t����b�2Zc���Ԏ�62850u�x�D<��~x����QDO���pY��y�ˇvN���@�F���QU1m�[:N�<�λn�����W�r���N�_��7m��%����ϰR"��fU�>�
��GȾT��%����+/ooo_�fج�a����@�(J��ʒ�NiD�ȃŇU�e�!E�6QǦ"���f��̐�l#���b�%J��X���#6�zX�ȑ5M[a�w�����,���Τ9����,��E9rq2s��	,H�L?���Ύζ6YTE�Kj�X�C&z��D��KM&�y���xgW'֠'����8T'G��d��`V�*��)n:�4��$��eY�'�{z:_�5��Wu�����xI�D��ux���ѥ��Q�1C�Y:��|���a��-���ӯw�+�,*-+ F��6�7��w��}~ؓ�x���t��+��4��k:�/���$�ܽ�=��� ��!��b�0dP�@]l�Q�F�����ڼ����悂�H?�9��lIi�i���޾����T�D�'��|���N�4��������S���X�T������3H�-��+
Rȧ�G���u���Ik�����c8����Bw�u�5�\��mWN��Dg
c�f&XXv띷�E3���HJ`%��m�0tMkYO�r,Ig��l�����O~2����$f�?޴=��-���������q�M7{��%-�w��_USZR�������w��{������N�tL���td�ɗ�P9�e5-}�e}���"�a�Z��y�[��	���1�ϟ�7�,)���R�����o�����Z���ܠRTVz��V|��G����K�c`�V7������cǞ{H�ј�0���׼�b0�S�����g�vl[��x*�ß�ۛo��Y��(/��޼�:�'-\x��p?��o޲�ZZ�<4���a�c��I>W<:��.++[�l��o�n��e�>���O�>�VP������F��:'�	�+w�׽-m��"�l�r���'q��:urQQ�ԄuX�@`u9>����^nn.`;�G*��@�b 8wG������L��W���v饗UWW�޹�s���d�ѡ���/�t��~��u#F~�{��>޲��^z5����Lp$+�|F:s�帴6{�i%�󲼂C<sM��K��O<v�8��H�$����?�NYqN����K.�?�\N�����?c �]}����Ν�QX�������H��
�:�u0'��q��5XNb�?֏����`����K�ߥ��v8両H#vK�����g�O0 $)��u���zӶDp�i���j��H���~�bv��4��{�9s��D<P0��u����I���8iBN^&p�ڲ�..�,�x8�(�<�a?Nsss__?��a+/��a~w�=U�5�a;��~Ӱ?���=���=��J�Q�c�UU� w����<��nkk���O'b�A�F� b�G�D����� `��`Y�e�4�d��L]smӕj�����"7�7���x���+��s�Y�vmcS=��L9�_�JM�h�Ħn�	��T<(;nBQai,��8�+�T?�3D�;���������&�t�ΏD#8@L���N7E"�d2�������#$��#|}H8]@��p�����[����7�nݺ7~��FOh�������:�bk�08� <X�ի�}��0[�G�6����+W^}�S�M�N	�A���p���b��k�À�x�iW�1����J\���W���W�$$r`��~���%����=z4�-`ګ��v����h4�I��L�K����Y��#ihR����H%"XW�׋�.?��/��88p}����ĒV��<x��Ν;'N�8a�DZG3��O�춦���;hHv�`8�<���ޘ�޾����{Ǐ��{/�)_���c&O.�(��Oj8���yp+��`yU�t��v�T���!��T���`gm��{��gO�2)K����.(�7R��1��zW�E�|Ǔ[������ude�t��M^�]*N��R��9�����B��L����S��+��@<���g�Z��J2��'� ��ŵu#������
���W�uÂ����-����^�� >�Mj7pJf���{+:�a��1.����FG��*�{Ƭ��PoO'V`+>��r�"�2�tpr������=����ȅ\�#��ԫ<���P@�6�S}PG�9<����9|��"˥X�������{?���B�8�I��p̌O�>��<gu�LE( ~,�����-��`嵁*�/
&�~��y��ʒ�缎�>����OGhh�ۦ�~��,�Z��2uI��fX�$�x>�g�18���r�C3��-�ۑS�*�4�~i)C���=w��eъ/+ί(����� �(S;L��XlIو��|����h��#�d׳����:�.���2|� �F�%QQx���/Y7(HlOW�==x��!`}9�Эߺ�ꫯ.+��m>�tW�����/���Ϭ3S�"y?��/3	�'���&��f����9�<i�Na�^��8VU�c�ȢE�탣F�Jk_0��׿��u��}�#G���7o����pґm(��c�=���Ϙ5���~%�.�e���G{4���S`J'��N�g	���s�]|�M�:�hZ(}����s��d�����o}���̲*�_�������ٵ�u
��j���x�j��kV�p�`�޽M� 1���>�u�U�p�=��H��C�pKD�t�8���p�u7�;�8�܇|�k^d=6�J�Z�~�Y�睡;��Z����KV:����C�7�;���e�$M�5�r���[�9�Ƕ��P2�@��h��f��
0�02;�����2�WZQs���=��j�Vq���gΞ1ߵ-����\Á}�(�q㦞�Hep$8�%��hni�'R� �M�6��+@l&$a&xj��!}�:�X@3��#������l"}��G 	��/xȚ���Z���ႂ�x"���Y^^5�zdcCӺu�sX$�z�*�38f&�%z�� C���C!��� �Ⴧx���(�����N����i#/6g,7��[w|8D���r�0�
����/��SK��jl8<jԨ��ʞ�.�%d�p,J�Ԧ�2�� 	((���@�,í�)YW���l=P�*����q,��u?5չ(-�xﾻ��3��,���e��قD_�`�+�*�D�f*�<��f���,�(4�wў�SK@0W]�r��g�.8q,m{��_y�յk_�F��[ƍ{�W���
QFňiSg���E��	�O޼m;�&vY8�XvFf^��ÓV�lE%Q���C�4������L ������}��XPUܹ�Sv��#"��x)�Z���=�+��	6ኟ��3�I�
c"uq��4]�
"��$J������:iF��+����q΅g���2��u�����p8v`Y���'=�x��d<�C��Y~߾�=��'�8=�:��5'��p�,�cB$�<�����1����@��Ҁs��+`�9�<�����'`Y�lq0��f7�wӵig&m��lF��l
���Ojn'��5U���zx->ůA����f$�(��13���-?�� �fY̈Gc�X��P��/*�͑��5�Q����B*ٱcgeU��3� �8^pTn�k���8�K��O�L���	��)�R8:Pe�(ٹ���yyy.���(�-x���^]VV
�r�8v��-��j߽k'����~8_�("}T �A�j��1+���� I��N9m��	��ɂ��^SSS*�3fLYy��[Z�?��@`3f�8���y_�/Ҁ�MC�O�mT"R�9�Ε����{g�;c�țo_u�7�ш����B߽@�S)�c��0C	[A���GgI9��	EyyW^u�	앮^�5.X���� �=�R��x`�p~0�kz*�خ�)Q�D���@W��:�k��@Q�UB�7PS���f���t$��SCi]K&��`x�EK�?�ܞގ��p6x�VS3nܸ�X԰L�,�L�,�k"-�`UYl/�d?_�⒎t �'��^,�R$)��9cޜ믻jڴ)$g*�3Q�#ŅU��3ZJV%�E�8�p{�<����Go�S�����־���|��*y-_�|�u��](��1O� ���nx�X4 ��+�=r,�/N�tT�"���\-{� ʑ� .�)r��s�>}δ�3���-�7�ܵ-�HT��u��Q7�rR�mo����n��C~�S���ɰ�hO��q>��bO�B Rq+��Jf���f�Y��Lxf	��}#��|
���#TVW��ᆰ?'�EasQ[]3l��&I��>>������&���C��O�����<��#6�=AF�7�F&�!gݲ��+.�t��g���o��?��/��Ξ;{�W������@0�@���~�����O>����
�,�I��d��>ڳ����ζ~)��e�AQP�XаaU7�x��Z�2}j�r�����{��ۆ�{�y�/��r��6�����ͭo��:�)˵?X��Y�9������s��;��С��)�>�h����3g��9s��޶}�?_��(�-��� 'O��c��=��3�ػ�l�����k�/B@��Ν7u�T BC�tm�?l��,�z�4etTd��%����͛ǐ.8�;v젎0�e ��uCWd��9>E�1Q=c�<�S��H������q��3�?ಀ��h� DZ��Џ��D"��$�[n���96@a��}�k�q[�`��1�өo0��m���@C��������s�AV�^�J';M�=�Ɓ��J�a��l����R;vn�s�y��a@�p����b��Þ=�\����9X'9��Ϟ����C�V�	^.�|���{���X�^\ZdZ��O?-*,Q��P�/�$�`n�̈o����z,97W-J�c�(\z�����ͽ�����EЖ��	bi���L�ܵ 򹹁��fM�2�!79|��s�njS���)������eڴij��ʫ�?��C{�焀��]5c�tx~�
�ܸ	99y�m-���ƃ\�X�O���w��$���b
���X��Iu�&M"2�(�����?��/6o�Dӵ����λ���M.c]w�u@��Zv;<f4��	��:���;��3i"l(�Xצ���-�-�?�eۉ龢��9ay��̺ 	,r� d��_e	��s�Hґ�Amb�k�mg���nw�n�����>�%�����巤��"�1��冂�D.���/��/~^RU��JY[�n��Ѧ-[��$#�;Y��!\v�)�U82���O�#��PnS�����T��u82+�l0��$$K��zhO^Vxzr�NJR��)�!�D���/��ٮ_��Ν>~܈�7m�裏���NK������,���X���[2�I�y۴�XNr/@M`���O�0�cG"S�c��)��ߴއ's���SVV?��mmm1-wĈ�ѣG3d�%@;L�Y���@vدW3����3�3 ���_�zNN��W_~�w�����:��Kcǌ�:yJ[��d2NF�Xt6��p����B9Q*W��v���<1�i�w ������
��s���t��֭---�]vYQq�C�2)��{F*��bF��Y�=���.�1m��O[O�>V	����y`����9B�xR�m��vlN&p :���V	,���ϝ1�@ XZZZ�Є���p``�}�p8@�R�Z�7ˎ��*�����x��[��Dc�c��!�E��0�m���)P���b�1���x�,s�a�e5���@ >��?���&R�)����� �t�6�ʂ$����8&�l��9kj0(Z�L{K��x �A���|�x�&�e+��g?+(��$�������.RŁĀ ��cp���
'�XW7���?��vwu=��Ӟ�ϝ7M�	�'�ZuÈ����� ����$�3 �*Dcz8'w���Ϟ��]�nsӡ���-��HЎ�Z��0<�R�Ns� ��Xpֽ��M]�0��p�=i�8x5�xDfUQ
x@'X�4���w�u��s��߮ٲ���4��OA%���'�� )���A����0L�n�XL���D�<~g��B�F���ͳ�e�dL�q�rs��e4�f���h�.��t�R���7�hb]�&Y�<{a �w,`�\2�ܴi�c3y��H_t���UI�0�}�7���X���lm�m���� ��=�����}�ZxA�\ﳍ�_J�R��$��5s�l	�ؘ}=��>�l���jky�>��]���w�M�{�u����>g͘JU���E�'O��K/e��`8�8����������h$7�(��&�(&����
_ [��uOg��
�P ���w�������^�WT[;BUd�����T���Ge`�N�@*[UO�BUU����A����
����~���S�X5��ڹ/�H�}~*(T3�./���O��w�<c�>GF�e1�W>O�� K@��A$\L��*..��d�
\
x����└��K��tZP䪪*��S�@3'�
v�&�E�V%iR�ad�3}w�m�>�>����6x���.�h��7l�g��6�`0Ǩ>("9>����l�)q��&o�c�8\i�Ț���zV3��X$����k��o��O�}����Z�
覷y�'<�H{{�i�/��x }>IYv��W^~m���t&,��/r�zYX0�U�	K��q5B�`]]g*c(��ј����Rh���+�9��/�y��k��klh��CjyU��Ҁ�,	��E!���2dO�@#�G�����g�A��oc;&�=J&8���JJʪ�k,��|A`z�?z;�xֲu�5$^8�|p맛�,=n��LZ������mz��_}��t"/��"G��h5��Ϧ�����`ǱK�$�&˂��
���'r�)5�r�V2�a�eK٤M��gy�Bá4f:���.�?������C�}Q��Q�%�P�D3t&/�,>��[o����2O�"�$������q�q��?�6!�ci�H[,�m߾�����r\QQ�>#���H���'�h )\ӡwK{ȹ��l�{�
-%�G�e�T^9��$�&H����CK�=c�5׮[���ܸa=2�0
@��
�q�IJR�fv�/�����y�Ҙ�%�YX�(�ۛ���>U4��%�Gԍ�4�KF��G���١u���`�׌�����%���? m�������++˧M��m��]�"peYҿH�gh���!BC��<4/�v)+��8qb^^^@U�mvtt�孭Q=��q�ݻ��޽��������|��fJ1h�E��T����⼱#J�xo����SXTp��_۳��f�$pD�`3�V�"��hqXA�E���S�̳^x��m�n���k�ds���v� ���C��C�bS�9�qRX)J�}I��&-��ph�P�K
�Ƣ�i8�SG�W�A(��N&�R`����X�����+oK�OKd�{k�D
}�(��7>�ERx�x�/�}U�k/--.ٸaK{[#X�D"�%?�s9`��L�U<�Ӎ����~��e��|*i�
�F��>Umm��뎆r�.���*	�n۳��;*FJ�ؓ��m{�����ՖQ5�n��I�Iwo�,�UP��T�%����r��8����˟oܺ���h�r?㙎����>��1b�5�����8��U�F��o����������	3C��ۿ��~7�Җ+I>pٚ��G�/�:�>��2�X,� l���QU[��%
�8�0��Iu��0BB��1"_kUVU䅱�ͳ�� ��?&��2�l���"��aQ5�$W�yFi>�����3��H�	l'7'�����o��U�����O7o7�N��(�m�7����V�qXR���K��H��89�ıp.�D,	؎�$4Q���~��b<�e<��F�����S�^I|��*w
�ִ��k�$�g�7���wa�*�\1X�i�`��N	͙��Aw�O���5.�Ȁ��D=�Lg˄���$�E�_���R�u�S;|<�(��D�@XX?�sJ~���Ǡ��Nk�Zw��6�����0����l7�1�l`8MX�B(
��SG�R�@`��Y��s$��hɰ-8�uaɴ��(��#(��#/ ��U�W���;�s�y6��D���l	�I�tHH��aWel�W}*�T2��t���;��t���g~�eD�]�|��E]�/��������k�|w�������?h�nc�O���w�z�Ư������y��pY��n�����!X������~:���K: >��j[p�Ȥu���k)}~,�b��<�D�Ҙs�lôӺ��5>̉Ģ��e���fF%�;`7��I�O��z�%#���i�F��b�8ZJ�Q����J"�ր(���)
8ڲ0?���˧�C�N3m��.����%�Ğx��>�[>�}st�$ԟ%B�����%EC��n�j̏Td)y�ۤ��؁�bvg�@8�z�A�`�M}ݵW]z��<�{����!MOO�>�vee%ϋ/��v���J��o���ӧ��@8�כ����+� ��	udJ39)ΩmZ�=�~$QSU�h4ZV�TT�Ez�,�C�#34�(�Y�H��8�5)u���*�5q�q[�j���������e:���B�đ�yy�睳���������A8�(��Z�H�瘬�a��]�0��%�D`�Z`����ɔ?�8��#?�#}]C����pEYuqq�g�?o�bx�<5�S۰mGVd�8_!��c��L����T����U�V��jn9x�`#|U��>y�QS&Ml9|(�Lp�g#Rjz�v�l��WC���E6�E�HH�	
kkk���eE)�nٲ%�L��� �EZ7���=��@ ��3d�r��:�g�8����d�	�bq /1eJ��O�������#G�-��K��2,nx[�h���z�e|�仓[Xp�^��E��w׽OX�LbDMj^���I&��\�>�<@�������N�z�����7�S��U��X�0����mqt���[���eg8�3-�O�	�QcF�s�M�?|�}x@��RyI��	l�G�T�i��[v��5}���_\ی��y����=U�Q��X<2B��xN6�֕+/"����N�-��ť��~�a6m���?=��ӽ��%��� GBU����}���Xl�}��䤃��Ɠ����bZK,[z�q�l0LI��RMnq�P�s�����7z�Xs�%3�\���2��E�VC���k���5�U�GT���$@�j��۷��8��e/�tG�0�]����q��,Y����������sXj(ēiɯ:��P<Gk&��������:}Z:c0�SS[z悙���a&�?���2 $���_�������6n̘	��B�P�`�����9�ҼAe�2E��s6`������3� ��w�5����$Mp����C��۷�0S��o�7_���E���<�?���ۗBU=Cx֠�U#��/�p�����UZ�@O(bMVT��`�)�<� z���.2�x���+��� xB -��d�!5�O�OQ0��&�-b���'�I�Sg����!�Ǹ�d���ܡM��vtuj>��xQ���7B[\ ���7�*f���W��(�`hϞ=�� #
���+�/D�O$�y^�J]��?����a�ĳIt<��F�����[���"C˙��t�IN*M��L.�k��0ibaQ���-����,����l<���� �,<eŗ�O�e�Yx:-���ې�]���d� ~^��h�Q�7xv^p�jé/C����2QI�DI�z�4��x,y(���Own߆�֬��k��1���V�����e�o���<���[6���k�gL�����k�aӆo8)D�7�Z����^�A	r?��B�I$�1o�y��;���h) <*��3���\,I�b�Ee��$�q�8��Xv����/⇘D�&чS��~}�@$�H�`K.�HU��@(��߅g@-K�E�Z\XlY:p�P�����_~	^��3pXEŢM:�+۲uT	���|�1��6�x���9R�5h���Q2G��g��躁e�Q\Xpםw���J��X�w��W���BcǎV�|@����7�|KwgWE�p�V,��}�����a { ��g�L~�N<��U�,�c�@�_I~��h)z� ���⃃��#S�*�w,�1$B���Q#��1��Aj�M���7�z3�L0(�eFK'|���'�"d;��eZ�t�C�c��N�'r��J��'�с|�{�<ܪ���������a�T�r ���ӊ�
�h��e�#C{�@M�\þH�?�2�LF�V�X��vضuxF0ªQ[5o޼���7�yDʇs&�/�z����r��Z�+--?~|qI��HZ2}��pkkkE尲�2��Xi"=z4�6�

�d����ԓ�Y#�@ߓ%�d�,�׍��̙�v��׸�8|e8�j���^�'�����^��U ���,��4f섪a��a*�ZUV��W<e��K��n8C`QZGK�o�������C�ȕ���vm2� �@�c���8Qpq̹E�
щ]�����M-j*�_׬` O�(���
Tͧ
�fM�6n��3

�צ��(] p�x|�֭�l��xS�-��zX���z�����D��C����G�i^��g�p��jx���-7/ϵ�z��G���U��&Vc������d��X(E,��E���}�Ǣ$�3Bzw���`{{'\�������S�W��kb��? ��u0����T4���3�<��H;؉K�ىP�Q�M�� >x����b���̋�@�Ȗ��2�L���ݲ���k�vɢ��OM�t��%%�=��Ԥ9fΛe���34#��#��%ն�@J�k�oz��wG�'�2Ú����KWn��t.9v� �)8pp�����JPg��Ç���]��_��g���{�Y6	7��|�Ft�=g@�ͤ2�[ւ��9����7^MK%��b�8ف�4WWUڎ�{�.*���I�����o�޳}��� <��λm�,*M��N�B�l�֗��d�')��"��}XVY�Spx{��h>Ԁ]�(�޹+K��Ax�֍7��=&o�=�������;w��ɬ'>��cYC�>�Ɗ��`A,S�c�S�`tMZ��ҒW��j���?���I�*���޽s���@��:�=;v�������1�>�( [�n7nLG3 �*�J��<y���c06ð���'�`�$�T�Myy9��8Y�d���4B��5�St����N�o�χñcǎ5j�����ŵ��.���Q��`�(�Z�`�8"}���̬^��W�{�ڻpÍ�5$-�f ,)w<������q_䉺)�G�W���"�3�++�QjL3������?� �H@�DN�O�eRL{KKwW�a#��65"��r����v�� �� Z%N� ��e.K�q�((X��*/ؖS&O��l;n��Y��` �{߉�)��	N�2�ȥp�*G	Ҁʺ�]42�t�M�dI����.<,��(
M'Z������؎9hy���]�D�� ���Q|2P>��@(D�כo��ԓ�K�Sp=xˡP�v:���#Q� ��� ٣���#�#��%��Q���nZ��|/b�}�*�J�`�)�t���`~�%c����}��\^������G��/}󛷱�����|b54�2�=��P�e�āb��Q�A�PPP ��{����l�E�ͱ������L��-��f��
g���f=T !��9^K�e	(z�N��!�����⡺?�v����oquDT�����QZP4�!|�2�A"l<��xqksی3��bĄ<+vm�[ʆ\��]3�R��Kt�8EU�F�����G�
�:v�ȩS�8���Ϫ��t|��q�M�b��J���� C o��=���SPP4r��ܼ�t2�z�ٵ�	&�ȤdvP�uT 2�_ы���l=Rm�͊(�����HU#�Խ����I��sf�|����ggU�UE�J�A��ȃk�>_?�XlOw,���;}ANIٔ�SfM�h� �i�8 ������iS�rB�tlߞ=�SO�o���g�"��hG�rR
���c5*af.�3I���9������,��\�`�9�,���åY�+�y!�w�4��fV�T��P������#�)+<����]Ј�yp�K�,��7��Tz&���G���N�|z`TI�0�d�6jw
؝��Py�4`9]�C8�����/��y�R"'���>� �L0T%4�Mbᢈ�aE��r�t�������e2�t�h�DW���3�]N�˲}ِ�@o��|�G����fc���`����c�aQ�ry��t����w@8(.^|n���/��fϾvX��\n�@�D.v�3�T,h��f��_�9�Y�&3|`���`��:7n�8�sE����'_}�5��Fj���g.�O������=��O������>���%�|���<��w֭\����(�Y ��>сOM&�zP!�a*����{�oQ ��V@�iv����M�I/�aXǉ��R"�Rq6,�C�ho��ח.��P达n�?T���{��u�r��o��[�|��_"g�pZ���lnn�'9.2W���̕M���}���㪮��^}�`��g�J
$��P��w?��l�G S{�s8��Y���]�ve(J:d���� �IZLY����������>c������+]]]S�NQ7��l���7�t��D��n԰a�(�3��c�mܸ���r�}�x�K�L�ػw�s�=w����aII�u�]�?�ɗ\r�$*R����_����nڴ�`�`Mh�P{{�3�<P�%�eե��:=>���y	Y��C�z���c~^�Fܗg지2y�B`�q@/Z�-�����P�(��ݹ}WG[{aQIGGOoo�_�4-��F���;���]{{{{�+���)x$���R=a��ư.�D���� ��Ztp��	?�`ooOYyɈQ#a�R��Oe%I9����D"-.Οu�T�a��4� �j� Z�4�1�Z��*A��Q=R�Ij)��,�?���x ���S^�T�KI<Cb���9�*�>�z��t�m�6����H.4�z`�p�
U��+��̡�N�Pq\{y��>S�ӚEn�8��T��b�	 ^��K�m�+%5S�L�Y&�Lc��2�A(��4���fϘ�ۓ������3k֌g��׷�zGyx隖dϲGFK���)�t���2��S8HG&�����`���%��"�G�/�ֵR"4���Jb���\G��Grk��L�L&���(��TBO��`PO�!�����ЭKn ��$`1Mv��P�Ab-�PQ�R�"��s9��ؤ �~~^ ?�w)܃��9}FEE�(�mF�1�
��*f1_ii�P�I��p���O���	��ʒ�u���v��ѣF��~�	6�\�xG�+&BG�ƑF.` �ŋ����!�M,��pu�e%9��T�Λ!� |U�@�(�G��.ҩ:�q���9<�3�!M7��0}Ƅ�P�c�	�ǂ]Hh	�h>�
�D����G���Z6���s��-(�fڬ��3yRU]M$O�u#c�I�P�~���8�LD�m����*�/������0P �B�i��F�yG�8h�"{T�%�\Y�+/��/��o�2���)�fȒ:a��PN~<��+
X�4S�LHKEeY '7�һ#��>�8yd�P�$��t�RT����"��W�b�yٲ�ﾢ�\���ă������lu���+l���@�JDvO�C�$�3,��|�~z
�Q�4P��Q��Pc3�Ep	��3I�a��c{��c���U�X4�	E�/��Z_�m-��"ژW�����jXK{<��k�k)pƹ�y�M��\�����.��l��C�����/�~��Z���ߗҭ�� �ˬ�K�a`[�!�᮶~�����_uӔ�s`o��)��%�Oa���ƿ>��=w��+����$�����˗8�������;::H��j���zC4��C6`����� ��,�DO��:OO���<�,�$����%,�㌖k���^ۻ�{��/x�\L�^�`X@Z�ETB� �
#�h4y�{:Ǌ'�s���O����nMhi�-7�Ruu�9��������Tn�H8��6o��k޸���fg+f�6��[a[8��T�x�����l�e�,�Ŝ�LIJ�₊��B��
��d�("�(���s)�L:�e��]��_<�X��fr�E�\X(�+�r&���,�ą�����MH����@|5�Da����ֳJ�³���G?���+u�x��ٵ�������.��o��w������Xu�i�ͤff���;����o.}�%0wX`AL��R����U%1�原D��ۀ����z$�����I��?|��o��ͥP�ptl��;n;|��$�0�W]q�>����zaA9��g>s��Q~X�E�� Λ�r%k��}��}�s�K���|�;1v���-[�l۶���U���~���W�H���_��_o۶�{�A����o�q��(�|�ry�׉M-N������
Ǣ�(�e^a�a5�%�I����ax&�gI*�'��tu�i����]������`I��<��ú�X����}3�"�d;^.�i'�!�5������D������q>�p JLd���� �	&�-��~�5�a����*2��f5]/����j��y˖�C�3�-��W��IlI5-`�6�
4?Q�
��В�>��.Λ�ԭ�농6/6l����L{k�Aiv�ڷ~V;�+n-�����iݹ�����#ǎ5/`aAǎ�%�l�]�
�I-
��仸��/�#Lp� ��o8>|���+:�˘߹��.<���."9�ʏ�~��0 ��_��/����9r����J@陯�'A���n�-�0�H,B&�	��LP�W+��Ш��n�,�*"�S��qun�����@'�!�FM�����^��ץ^�V��$E,X�m��I���,��G�B9.��Jbd��<ӄS��2U
EI������{��+���٣nkm���7��Y�Դl���V�,��>�<�4YҠ=���L>x��8����6�h�U�͛7�y~o�Tb$�[�0:�D���my"�������ڙ�ES�H�T�0��L��ȡC��mܰ�Pl	@�Y���{���(Hgm�D5�Ma�H4�`�E�>�/�[�;���>���L�c����[J5��eǭ˺0;W"E��P��c�2� '���� ML����\��vjz�ر���	^��\l*F���%����u�=�����}��P��G{������h�^S�� 
�xg�h,S��]�
ײ�?'J�X8�&&gAT�}�\y��~��}��߶ݎ��eM�V���h�V5�ֵ��t�����<����~lɭ�6��Ｉf��3Ŗ�\�|��Q*A��L4�Q/����e�����`AOS��g_���o	f+�Tfrl������a=��_��tQ�yn�2�.L��X,��q+�$!:�*���'�1)�,��6���Man
cҾ��~(C�Gf� �F�N�ZV��3�_�K�6�Ѣ�R��Q�|970�����T�(�%9�*"8�Rad�JJ896��O��C�{���c[[� �^���:�5�� ��d�����*V���	�Ǒkt�x���~���m��w����t��2)�R��ݽ��_�_��W��;;֌���H�����
�;���'?98x���ոT�9�V�����B[)��j�2-�m������o~��c�o��O����{ld���C�����w�9�����ڵ�s��@�T]��E����Óp�
��#~u�4E�?�o����xM�^������}`׏�����O��o2�Φɩ���@�
��k^s1�~!�I����������oq�;�ݜ�q�����<��<6Է��vݷ���>���w���}}�&Ƨ::�}���ۃc|zf��o������5�p���3O�z뷀0,��bЉ�q���n�e�Q���|�K_*
��3���m��:g0 ؈�S���n���?�K'�,�����\w-ߧ?��}�3���h�7����pe��kT2�'O?�����_z{{.��R,������!]���O|��{�1�r.��ؿ��K^��g`�[n�ڧ?�i��*Cu���y�D����������M�W����'Ԁ�n����w������pÛ?��/`�2C���|�u�>j� �A��]�;��suʹLcس����}tF@�PgSe��Ca�\�T�8�������S0L@��;����z�����if��Od H��U�E��@�ΰʭ�� N5�n�9ۦ�-�A����
)�,H��W���V��O�rM��>�7ܪʖm[��c��V6�14ժQjq�����-�*l��Z-����W��w�s���X��<��_��=�������p˲��s2 �d��'9�3.�XL��L]�t���ǲ��?|ߣ�y +��j�
X"�i����c�<�L��^��}�'��E�/����׆��Y��'Iz�h*!��f�^�c�)ad���*\��;uǮO��pR�I.�,5���^�M��$�-Ѿ�<�	�I������T����Ż"�2��Q���EA`5�=���t�7�o���&IG:�
��e���	a�S���V 6�D7u�Vd|��a����gM#U�m˷��{n����a�4�Q���-Q��F6�Y�CI����*�s��[)���/pB��C��������5�rE��%��Oޡ�l!���:X��k{p�ܰ5�_�w=�a��.w߶��%��]�l�g'��e/�W˙L>��_v�eC�G�;�o?����Ҷ��3{��i]Q���1��}R�w��k�Ps5ɧ H�[����O=�d��'�o跪s�t�u���^b�m���"������#����S��㲒���1e�����S'*�Ņ�;[��-����cM���l�jMI��mo���|S����f<���GaV:;���e�����S<
t��Ï_��L&�����w�����>��s��0ッ��2Ux� �}\��t�8�V;:ڮz��n��O<�2�,����m�S���Z��fەz�Z��)ͪ�
�傆�Ol����I�|����|�6���b��4&KΤ��d�"�`�qӺ�e4S�t]����w����+r�m���n%C7�R�&�Ʃ�h�3(�#>0p�曾>1Y�d�׮鞞������|�ۏ<�H�Jppdd�N�����k��O<q��a��W��"ZK֔��[Y_��>��矃Ca������a}����W\s�eWq[���<��A.���������o�֛�$��w�>�4\�g�U����e�����hkٱ��n��x��W���c�����k�+F�Ǐ�q�] ؀ ���󖷼�_Ͼ}���.�-!��Vn>�r&o@�t�g�<��o�����y{{k$׽�-W�ᷲ��a�(e����}�c<>��ڊ�y���q��7����D�|�-����ej�$x�G*��%z��~�������?�fM�X�������G?�O?��� ��"����6lx�k_�o߾O}�S>��i��%�������a�����pa��|��n��V��[�u<x���o����cĦ��10�\7�e;e_�N��ɩ;�c۶m��$o�{��~��{�	�SMA6M�<���߻���������5-�#c��Q�1�0�����xH�O��g�
,$�2w�?44t�m���u.����ȸ6��G5� nJ���R^�j���2�F���|?m�ج��\�WQ݂Y޺u+�()��CQU/�AVOe3<G�5�\�R�%Zo߶'����޽{��R/���S�,� *�`���خ�[|&�ɲ�C�<;���}��P�JmC�dHX��a����,��*��u�yb)���i�(�4��[���i:9֩;6�٬����Ɨe�x�B�,�DG�+�B��1�x�{R�����%*`})z+��`KKe8[T�녈��@Y�S,X!�|�e?�ܐ��]��'���+��\�D ��4 �U����?��.�Ő&����&�4A�6�^�!Q�d�2=5��:ձ�^pJK1�!��Y��]]]���ru�8��gJ�x"A��Ls�S6-39�Ո�<x����Tk[���:���,�$nOh�Y|9c['1A�X(�Pw@!�uS�l|]>z��C=Ң�::�/��1�-P��9��V��'B�(���J��q������{0�.�u��������B��-9�77[;�ض�
�[p��$8�T�TlB:0���48¹��D*:@6�ƣ*ԗ�����o��sv�S����G?���Aֻ�������-��3˲���c�:���֭�)�1r1��S�SG���b캮���ꊢ����?m-�_x�ŰH�m������x��s���1�^2�YQr��&��U�S�B�b���H&��6�ٍ�`�Dn��aK�VXu��~v�-:=3�kҪԈ]��Vu�@J)��FV�?(�O&�/�����.����c㡨�n�4�����T�K]��{�oll�OU+����C�G��)�Ȥ�?86t�M7�+>&IC�� ���\Wd��,]�3������֛͛fǟ��{q.�'[����ȗ��eN$`+��ַ^{�ss�B!744��/}���8*��~ٶԣ+��2��~���j�����[>�/�fSko�&���L�l}�S�|�W�',!X����{ǎ��~�|��߳giI)
/H�碜��

�>�l՛o�9�˽�]��P��}ˈ�z��?��/`40�`)<_��wq_����,"�� �1kJ��]���o���6o�ǋ�>k,�]e	�!����l����*x�=���A=����{p�~��x�g���7�ygg'��哟�$�	3��/�%F�_�"Fc��o�СC�.9�#��w"`�����}�K�/��}�s�j����8�5"B���P���z�;���\�R�E�z�'�Yjq�z�m��/o�Ϸ(�A)ߵR��O�&'�1�7oߴi���L�Rݹs'����w��<��@~������d:cb�����Q���� (45 ��g����`�yUXGG���(H2V��]�X��j�@�q"ЊDNF���t��J�M�x}�tl��~����޽�xO�BtբC�I���1Y����P���Gh�
"H�U��&j�7��DSk�B�� �5�@�	bi�5�>�;_���R&� ��忢�a`;u3���g���K_���i�#���ͅ"� ��"�[Td
a$SW 4�ᕎ��i�"aלE��U������X�BQ��c0AE��oK���'D��hK���_��P���v�Z�̱�c��\x�]t�ǴB���\���Y�}*������c:��8�����: �1�@�+O�i�T�fD(\���2$�$�U.K��4����������/z��,�X�EJ�����������^P��K���rY�
�! ����$�4P�SDr�0�f�^�N�� ��\f��5ÓSu��[���Ǝ�6Q�uEq�]�ص���hJS/�������'�<�K�xD(�j�C9�a�KV��)��,���ۢ���FY����v+�j�?����ă#��B��Λ��a�`�QhU�G|⑇+�r1W���+~ 3(�4:2���ۓ�g+�3T�tB�L�?[�Vn��m�����;6I�|����Tke�&UY���]�JC�z�b�@�f����E����_RC��@҉]���Eeϰ�ǲ%
�l�\U�+��Pl]��v>�]^����t�o�����g�9L�������}��,*���3�2c���>QA�k�����r\N���|n�C�k�77P�8Q�j�9�K�tT�kPPٲ@��=Ͻ��g��M}O%o��׭JD_��?��ρ�
EF6���u�q�a<p�������3�@K��`���U~�[߁����>�yS�mWҙ|����NO���g������Îg���?��O|�GS؃�_�����[��$SՄC��|�_����y�~۶m�ѓ���?��]w���'��M�L��@$����O���[����;��)+	8H�}O(�yP���^��o���Gy��������<����Ph���R�2T}�T�y��aN�Hy�ђ�����?~�ĈH�����x<
O���?�8���t�PēUx���
Gg���l���[�n�z�UW�Q���|�����o�?��P�ML�ג����J����?�]�a|r���glb�_��_�`��
�����`PL�r�k5|��ʹ`R� ���eG���0�����d3�s B7n��NLL����$���o܌u[�W&&���~��},�H+�熆=�Q��9�C��s�;.IӔ_�����G��޿<�ܝCC0�k��vwt������\C���3sG�t۾}��@?��O?���6��:��}T�����f�(��(0\�l�Ƴ��,x>����L7�x!���ҜF��JRm�ɦ�-m�L�s���p뗨�	'��r�o,9���pP�ox�5�\#e;d������%EM�?S�#Ir/d���Y�h�>��٩�T[K�>�U�������0 ��>��r=�.�r	}��#��&��Ia����B���r��fޑ��hH� Ự)�9�I��7�O��I�+R�B%��LײB�^(�R&�tq"`X i-�:�e2괧�����S?[�Y?��Ը�E캾Ȏ�����b�L����� HA*�������z��]�.��/�AWvҟ��1�}@��$��C��*�*�6� ����T�@�q��+Gq�D΂Y������z�z��tf���-���j�[�y��(*���ޒ�vvT��[�{��s�ݑo�y��/q��u|��8�pP���\����,���bi����ul|��/���9�sλ�O���3�`��ر��`�i��zK��T)oXߣJ��3s`J�����]l����zF׍�.�_�N�����ib�IZT7gfg~��`����?ٵk�f��x�o����t��om d���/��2����Vc�Kg@������|��hfKq{�S�#t��dQ�r��\1U��K��t��:�n@Ev�P04�T�j���䰢���_��G��:Tt���M7�߰)���*�v�(?�B�A5=��7��Î�J�U�q�n�0CG�f0�.��f���Ӆ�>�*��'��4.7�S
5NcIW>���~��~�kǎ]�lKg���=������ X�Kۆ��{���|��rǝw�Pd@6b|cղP��q����S�cY�|���w��w- M�m�׿z Ԃ�e����G��z����b	�A�teII��]�L�׀-�z��ћ�r���{zz*��qދ��GD�а准��u g�ˁB"p��[����2�i�9�oy�'���gSohޖ�P�����P��b��t�������	�p(�/�Z���7{��g	c������\�nIݭ�5"E����ݻ���?���}��o~3f���Ѱ>�.����Z�a	n���$���k����s�!K�V��Ng@G�o}&�EJ�����iv?�	hNԟ�a�D�0�4k<P�⹡�w3�����pO���C"U*�o������������#�6m:�k>�.���v��߳��������:X7��.��s�ݲe�$�[��6Y�ᖖ�r�rx[���G*�]'tl�E�!�G-Ea�<�g�t�|>��c��r����cD((���K��
E�����#s���^�M�Qb�����~��L�۞AD����5�j�EeR�o_�<��az�{��q*�b�+��04��IRsC�q���g�E��yR�*֮Ï�D���ӲcNE�"�_���;�~���T�Y����v�T3E��(2�v��,$J8, m
06�\�����g���+7"���+
r&CX���u����["F$�C��X���Itx���
!BQ�%�+�������#�29�<877�rZlN�9�w}Jv����0�.�Ͷtlݲ��K>%��������U)f�/RiٲJ��fә�������b�%����l>��B%�_�t|�x�+������'r�D�����'��N����������~�o�;wlJ�i:Qd2(�\~n��:���º�n�ך�w�NN�+��틟��mo����~�\6�^��K\F9' +^���fo��ۚ��Rv�y�~�׼�s�t�@�Z����~�Ş @�z�nf�L.���<�����&~p�m���3�|�;W惾��CNʼԉ�vm�hj��nر��@�\�����ӺXli�*�*���������^Ak�����-����LOO���뜱{���8a�Rd��#d��RŅ��s�N��ݭq�T⾷�����wz��H��P��+O=����>���Llh���ܬa�Ȥ��aXX�~��w�����ue���^qd���zF&R������h��9><#����������豣���&^���rI�T<O�ӥ���>�OضL����\��Ջ��)=\�c2�V�R�'�1��Ⱥ~p��AJ��t� f�<G�0�aO0n�Z�CL0F�X�Eɋ�I,������}�q!�r �*y#�h�@�XJy72��x��i��#7�c^�)�W�H#s���2C�V*al0���X̯�W���ށ�?�OLMM]w�u@��>�,�c�p�jX�}y�U��~����=�B��_����lj�U�bH�bv���d�ŘӶ\)۶�/d�����:����c�S�41|/^�y'0}m"`�[��X1�3M��>rs�,���x3�C�h��q�%K�;\�?��޽�,'x��Ǿ�AE��J����ì3��P�� ��������޼ys�2"�E�w�x |�-�(�n����f2�B�?�}��8��'J@���"xՊ �-9�ca�6?K��s��Y � s�
��jVC��eQf�(ȣ1ej�x�J�d��F=oUE�TK�r�G�h��,ܷ�~i�5���qdT+�0f���H�4"D`�����F��6wͰ�)R�#���)���8w���8��Tߺ�⵽=B$)��Bmƍ90�W�����D-"�9�֭���C�3M�M�il[q������rj\s�	�0���$�N��U�T�˕��Z����Zr���l.��#_�,������A�6F[�\��\��o׮��>p�����.��_ H"���\�I�$�ʉ�	�D��]]k��U�qd uvvj�4;Y��7��K�&
jk���ږ+� 029�{m/����4���8Ui4�d�(n�������!!�mZ߉���ֆ������Q�^pqyE�әT�X�fs�@�����<����@___�
�������F���%�͖ʳ?��O3���6o_S,�	�`��P���f����q}�`���Gհ*��c�?��'O��	9�YU�$-@.iMVg��������-׬[�FVB-��Y�v����ѻ����W_�ۿs-τ�-������s�6==�F�$7'kg|!q���h.�,	������gS�jQ��)Y�l�rH/ya>��G�S�����h�k-Rv������`���)3]��(+�畱��������R��,�����j�H�T(�C`���UMVDˮaGd��I>Ų$�03eX,k�oU~����������fO�
I�H�m�ژ⇇�q\���Q��o�Q ^��+=�o���0]2���O������/�6�RѮa,��snÐ �iR�0r�w��f����<%���i�G�H�����y8v�PrW\��a�
�U�m/�#�V������:g������ْ"�\���)��9��wXvXlk����$Cx.��|6y���ҬQ/��;33��D��?R�y�*�8a$َ,�͙�h5�2�{h:�E�-�nUY�VX,�w����<����y�6���h(J.[����`j|?<7,�4u'��m2���3��s� ��Wx�@&lp:x��X�$�q��k�#3��(/�1[%J��V��691����%���HӒXs��9G�EmU����#kIb��l}�s��E�Cx".� �yX�dZ(�!�)~�	�\_rO7<M\+���)Qj�OJ���F* �ˣ��C��&�b"%�S��]�A��B��,��NV5G֚�trrZ�;����K0j��K(8«�,ɚ�+�u����X0���酠��\��=x��W(:Q�{�`8�X�h��6c�6�B�T�gF�/�,{��A�HB�q�\��ƾ�aC��7=Y��ݻ����[�]��T���O�/�ix/�����{b_`�yS!�Pq��XQ�i%�Me�\6ֵ� �^&ۢ^�b�b;��m�\��ιj%�/
�GuY����GJ2�I�(�k��pH�Y�أ?��S����ә��NqIG�4�0Ru���=�O��ٶ�v��e�9�q�v��r~ӦM>U��ҚR(�I?�ө|�n1G����7�79j���ι�� �rl'�M��)�N-WWUR_����&i�=64||l��w���Ӊ��\2tz���{���W����V�.K�'+��k�w����et-+D��´�x3L�p�G>��3ӹb�AI��B�3�B�oaPr\�L�S��%Uҽ �P�!���X�$
�3�/��2�,�-��R����/��EE�fF�t��	�#)�*�5i�J����1��#Q� Օ���Ӯj$D�:��8�fH��P!��N��8��|�
o�J�ǭ���8}=��AꋀJ�0Xl&�۪���w�9U`�F�RƸ��K�Y�-�rxwN�`�)��t�Z��j��!�5����qI%�4L��8�8����pZ��'�۴R)�w�`��[(����ę���*�A�s؃�*��T'�b-�%12�-%J�	j��j�99�X߹Igzz�3��L&]����1A�橕�����1PKj����=�!�%0S I7��ıF�ac9Q�(�ْYN��C�-U%�O�&���?;�g;u����9'��0u]���%���Xa�)-��nS��os����Er����s_��,0���؎�+i#�ڼF7��Bvbr; ��~&C�w|�s���œX�y�8�?� g	&7�g.*����,%l3Eri�=�:��M�Zay�-�k�E��H3qr�p.�N�ł��䂛��	��$] ð����ly��݇�t^;+2�� �Cْ��ʁ�!�|#���鰱IL����nrO5K(b��q�T@�{���T������ӓ��*�2]XP 4�����pEJ��2i8US����H��@�Q�$G��Ĝ�:H"���e�UܾgJ��1A�C&���0P�l6�����k2U�����:�5B��a�aeY3���fH֣�R���U�Rd
J�*?�Ԑ&�����-��;`"^� Q^�@�� U�(���#;�	�Z�0�k�w������m��slx.�� ���9�=MH��+Bݵ("���SV���]�ҷqXS��O�T0���Q�+�R���B��N�\�e򢙂1���i)f"Iٺ��b�U��:�Vrad}�"�|���k)��UX���-c���j�<�j�f�*3Ů�߾����kG��b��Z�@�o�eK����z�|��B�$����m�B��c͛�֩fq�6z���|dͺ���\%�@���4�V�i1�Pϵ'��|��/���߾};�ă����`bοb�,������=��À�\���z$DQx��+��q^q1䢣ۏ#Bm��<��SKy7�00O��)==
�ss��{����i��O����/k�։���fE��Z�j�,�OM|����'>E!rY�Ζ�<������kw�e$�ީE���;��U:�-���_o|�ߗ����|�߿�Hd�W���(��w6hy��L��5Z9%��	]�*\D����Ĭi���H��O��?�1\ITL��?Wv�q�E4�t�:cX!�"�	�V�T�K�
���vק�a
�I�:�� ^��_`�� j�����s�)�'ӳ�|�[N���:�/a�V���K�Jv�\��`�Uq�%h&�t���wq��?O
��<gr�-�6��� f�䛊D���ɵJ�:`g��H��� ����&Wl��]��}?��&�8��M�Ы���"�I�:0Ε'Y���4�Îm�̲�jf`��j)��-kq�:�6G ���[��zx�-�j�Ǖ���Z�d�2�t&���ܵ:�O�C�Ԣ�1:�ᓐ�S/��/{��T�$��5�P/e��L���2Đ� e�qH�$�[����L�\�T�a���aץ0Aȍ�c�rP���yA.ه����"�v���l�������׷Ĺ��C��/�UR�$v�YP'�ua��ȋ��k���0�f6Ήe*�G��Ĥ�$���^xᅁ��]����O��;[*� 	ˁ�E����QPȵm%s�B�(�r�uk�����<P��#��,,��q����TPZ|�WܾK,؝�)��*�&�����k���SO�I���ԣ (�=1�X�eZ��pa<�H-ˢ8�Z���jwg�wd�8����8_�EpʂwZ!-T�L`G�#3v�MR�j
_")�M�{C#��I�y��G@�5\��ͦ�TjϞ�#���;�߹)��DߝQ��֎��m�7l�e�'��8'H�"���>�m�5"�����~H�l�Ƶ�+����ÓSs�lq�J��YB����[�(������.�������>��`@`u]�-�Y(��yi�D��
C�GQߺ�7�ˊ��f���b�A��fj�j�ئ���ڄ�B+%���
�pl�鈡�
yen��/�l.������4k���Z�'�W����J6�� nܲ��/��]�),��ti||��~�����ᑡ����=��;:;����h�*�_x~��Ç���2+���9����Rl���j����1�\�F�*�%ef�,j����s��>B�_�"�ںj. 1jxÚ�\�A���|��屔`�;����C�&~����uc۶mv,�ݻw��:thff�4S���-������=�յo�^�r����-�	�����27��R� �M��jM�B�� ��_�r�����_tB�����2~�y��U�{I�G���fZx��=�O���]�J��Pr�k�4v�r�k���Cb�v�����Kx�_�%��g�}��b����U�۪'�,(H�%�YU|8��Ze�'h���B�:3����E�}q���Ƌ��_�#fE��H�܀�v�Wo��	G���t�.��K�KV�v7}Bp�KH��kx�`�e9\���c>ii�{Z���^N��K�I"�s�fgg���t���u�Ә�Д+�=�I�)I[`��Z����tU�D��׬Y��V�����۷_y�cS�###�<�.�$ȉ4Zv:�Js~��YY@��R�7���[����)����7-˚��[�)z�/OjSS.*�RYr@�����L5%�v�^�-�jF���߿y�f �L�$�L4oi"�&��&���r�rde����bYA�6111<3��(
_u�$��Q��XX�7n��δ��e�yA�3��pW�$Qd��U
!v���ӓ+�@(�jL(��k5�<[�})��F�ߢtbR�'�'��}�ַ�w2/���?184���e�X�1%���"��D�k?dY�bX'�>��$�tAWtٱ}E7Ͽ��L�ej�||l���A �g�}�ȑ#���Kg[�6ﺨ<7�����߳fM���_߷qs�P���ޯ��O>���^R׫�X��JuyM8,��$Q���$�!3�g�iN�iX�8Ҩ(�a��p�cs�"C����Ph��c��PsR
M���� �
4�W8�կ~V	K������¿�fR�b�mrr�T.1�����6ˊ1=\`��^��.�g�|1j��[��&��ݘGi�������G�O�(���`^�O�S:��I*�2�8,+oz���b�1�mD��F�qi�[^�ry�lp�%���hŗJ����JX#PI���(�of>q��_�q�����_�KI�y��՚��yw��/���y�"W?i~݊�*9�e��;(2�\���Z��K���O.���B�S���[fQH���i��Q����$4OQ�8M�!:��v��e�6!{'l�t����U��!�)�zN�p81�*U!�tŶ�P��-8'���s_IݗɁ��F�����$]M_4g~����������N�r�2�̦M����GGG�S�g�II�;9��e���ce��BZ� �0[l���#;��,�0������QI�l(�*Hb����i"��t�
p�����`Gҥ�� c�W���OOC}��P�H��+3x��F��u��SxVIOOO�t=_W���`GX��H�!�ngڸk���M�CHĶ��
Z�*o����"m���ٟ��>,ߑ���`�����믾��T�51v��?p�C�/tw����Ng���|������h�����sg��fAb#�fm��:�l'�%��C�%���_)ds�U��~08xl����al��Ǐ�b�tvi�z�����?~��?�������ٖ���B�����x��0�=W�5(Rժ3���Ry=p!���LD���PY�%(|YIL�	�乡.Q5��tId�?X�f��7�IS�|��|�Ġy�&����L�������4��N�����I�ډ�qQ�(��Dhكa9&%�1Z�$Wهg3�s�`�KR����ERSX)��v_@)59��f0��9a@�v���Zf�؃0OJ��1ucz�Z܈,_/b��x�r���U�.R�fINRn-�&1��7��:c�D��O:E��O�pۉ�4�I�����	��G,3�o�܇��z߻�b�hoa���]�G͖	G��t!)��:����=�q�����i��E$&�/ԥ-I�d���OfʈB�,{Sf�1�:�˵�5���63ө�E5l�$�r�I�(&�9�GHtBAL�&����;��Fcg�J%���(��\�ꅀ���H���X�V�D$� �pų����J�>�r�<���T���P��K�U���"
#���,�t����H�����U��i���<j^&Z�����ؽN�ü��:>:44������l�E�NUt&qh���Z��TJ��+�C�<[ϻ`��sݺU��1}�Wb
h��7u���F��q�j�B�V���uCVU�"lV�w!�}��x~rr���������K�����C��CC�ܿ��L�|#md���б�܌$��
)�Q�x����^$x>� �bm�*����ȡ`F�\����s���;333"H��I�D��w��{���{�a�Ⴧ0��c����ص��ى1ؓ\��ib|j�����yfe�KbxV@$�������0�c�#�Lp��'����'U�����
�j�X���ݤ��5?��xP��DyJ�GT�_/c�4U�dI#��:>Ѳ}��倓[*=�wRx�!�J���}Q��R�y��8I���Ԉ��>�X�M\�%�IM�_�q�����J�I��5]�|(�9�O�Wf+�;6�#��Pީ0�C��O��W��T��`6�6-�^M�%j����b���J/Ţ]�H�����>q�Ϗ[��̮�&:�GƐ � ~=��KQ.�F��Kl�Wh`ݼțC[�J��Uݐ�$���������d�v��u��	X���1M��I��tzB�	R�T3$1��s����}�G���9�IALO��\ip��H-?V���y�t�4%޼�p�%˚���I��I��ĩ��#��+�v2��wtu����R���Z����)V����dQ��=!H�)C0�Wx0�i��Ry�P�s���P��\�R.��iV���L��(�m˪s)$]���[I�C;;;���j�4.\w�+q
��������4(�,s��`Aʒ�ڭ����2��!���m6੃��\t)���{�7CG�C�K����ز��y��R(�SaÙ1�<��m?6��H#gC$�^D&K��5glt�%-K+Lƶ����Ȑ U�=MV���k��>�́^�T*�[��C$ٲ�u���OBa:�\����K"�{ְ;�� l>��/�MJ�����*�	ք��!1�$$6'^r
.<f�v�M��R�%�,�%�0-&^�+3�l��J�<��u��a:��6�((����|0Zf�6҈(kSx	Px��.�!Oɞ��g=n��jl�E��%]��?YP;��]�,�=��z�ǡ�+Ę��_.�Y}��v.�|@dA\�~ቝIz�4���Y�O2�ĈxJ����}��yP'z�O^���&�D�*$�J����tj�xѲd�U��*�V),.�)*�z�d��Y�fa�$����"r|��K�vbq`L�Ve�N~��-4��V����<�X.��H�2"!��<g�%!�|4�ֶ�jf�+�Cr��e��\����%�G�x瓊]����\�t�	r\%���7�|�0��uuu�"�B����5��4��^��J���i7D\[<᫔��#��i2�>늆WT
:���M��R"��g����Y�	�+�A�pR��̵���m��I��koo�M�N\+���F���".*��=d��R,����a9v������7��WGP�n�'��_��?����$�Ϗ��yI-��B_U�.�HF�w� �u+wd�8�	��J���:��"���z��l����Z�z`G\fQHt!C�q<��	3����q�B����V�J�DY�b ����Ɋ��*73�P��.��>k�
�Pb��n&�/�H�K6cQ���7�Y�}H��6%Q�eϕ���������^|��D�y��{\'d!�V��T�$�GW���%I���%N��]l:��T�U��r3��ø_��dI~����FL����?ᤌ��
'x�W��j9 �LP�g�hE��R��hi��~�׃U"B|�Eq��]\zq��h^�Ir��	�p^����W)�Ajg�������	5�e]�G��� �� ,��`UXG�D/�5����1�P#��Ϻ�
�f0��3s��ȕ�:����˫(�_ʱX�z����B�cu�?d�)�΢ۿ"q�y����մV� Ph��y�ļ�8=]�B�.R�h2�K�
�0
���\�ՠ�B¨c���U�Zn�*��丱k��d�D���zsh��d/A;����\�2�~�w�e�6�t)�P��uT-�QI�@�/�)L�;pؿ�5���(*0�˚�`��|R|���g �a&ϓ��J��aNC��Hk������������щ�����M4Բ"��j�g�	���j���x~㰏�=�'/�rk���oo'�ub��W0jl���;�s�5n�p蘿n���ҭ�gtv�P��S��I,��<*������S�W�&���˯�Rx�<�n�Y����d,�����b��e>\��>XC�8���Q�?r\��}ھl��hA�M�<�uQ�X@����Z�S/�0`�4�X#\���KWW'�<����h�N�aF@���&�K�Ҋ��+��׭ k�f{u|��IY����j�>5
�T��碦�i8�i�/���:��-�J��Jg.-��ѣG�_�R3�o�*�-Q���'
D��o��'�DMze��̈́�	X��φ�[�:'0W%](}�"P��\�O't$-�@��PE���Kp�y6VQ�Z�Ḁ+��gK��ŕl�S�/�|�rz,�(���CM�G_���)#J/��H^Ə��A�<_3QS������{���H���jr��W�%ϗ����ՊDHl�S�����W�4@]�)�ASG�#yFQ>����9b��e�E�N������dgX^5e��H�yy��)	L��>2 vX�#ބ��%�i#�nH�3T�pU�ZC0:_5.��R�P���w�CV�A�%��|C?3^�/a	���i.�k����a�z�zq0�iYH�*{�bP�Z�����IY�f���G ��r:�:<ϼ��LO��HHt�i�I+-�n�?or���C����L���B:��W��d�I� �v���q1L��jKd�Թ��l���xc҄��Z6
o�(6kN:%�/R���tZ�I���CU���)�IH�9�L�3�&�K�/ю�/@�pr��i�,Pc"O�*q����;=F�D��Z�ʹ�ԏ��^jd
�Ȗ$�E�����M�'�&c�Ke�R�0�===���9�8��a�p��Q�L��Y��uR���V�zC�O��Sgg;�\������ns=kvz�Z�x��$c�G���ƚ�!��ؠ�iB(k���Ro�(TJs�0���j*�o=�g��C���R8-��2N�v2RgC��T*#�)j�n�2�[E���l	��5� 
,):5�=����-� ���E&^���w��;�`�U�r�n�����MW�ơ6�QgG�wb�� j�%�bhk�%I��@Vӑo�G�Ϫ(b�Ni�g�2����2( '���nhnŚ����y��?Ʀ~��������s1�?+'rX��0�D��~J��	%�p|��}%��tU�e��b�$�"	����am�Z�]dJ���yɣ�孥FRM�O�e��8�U=�Pp f#�w��Y�B�"�����(������zqG�$����DvaLJ�9�b(�k[:���r�c��մD�>��i�EA�Mr��\��N��b�@�j������A�����ȱ�t8�H8��2�nv$qE~y��,�(�B6h�`'x~TQ6$U�B��Hb��>BU�"�U��l(�����@dSJE����BKH�d���"��W#Y��Əz�c�`�	�#k��	
�"��^���:���!���W�J>WJX~#��F�MW�\ZWU�.,�bASI�T1��c7��X�2oQ��[�n�	�\�#�XV,<�x��"� �)�4K��\�a�J��+�ߢ��kh��_��+�?�a7�}�����<���Q���WY�|��5�:�9���"���)r���4�m�x�#��	�Tʌ���<?�Z%����E��h�&S�ξH�S��F�P�i��C��Y_O�:��C�u,�sd6;a�S�n�z��_�>u�`v�4=;Y)�(r���Ғ/(�0�$���iN҈����������V(�rr�|�0#Yr}ofzҭ��[Η�@�\[��zy�<3y6vw����� ����?�')���3�,��<�F�9HF�N�^��H�����g5j�`+Σ����t�i�.C��-i
��aVT�Ð�����(K'���1����s@b����.m,s�)Z�)��8���$�So7j��R�("�-"Ңi�O�o�e8 �1w8Y��ø��<���R]pT��ߵ�q3)���WEjf�ҔfN��/V��Բ��;lz��V7R�|��fk>�x��X�|,fC�N�@}�Z�X'�\�5��caf29Y�at�NYyd��TR3�p��fx	C]�t��`�i��s��+��+Dx�N1j�+��B�"���	��ȼ"��F�a  �.�"7�o���^m�;�ϴ�h��V�X �e�=Ǳe�0�,cJkd��I���u䜐Cp��e����TU�)�.�̺g�T�D���ܴ��az5��I�Ϝ���@M�	�T��yY5��d1`�����T*��g�i�4�6����h�i�bG��%\���L�a��b�����΀�Ǽ0�"��0�-NP6l�a!�҈�(x�s��Z���d`�ZI�>����tvt��^�[��c3��B1���Ƀ��)�|�x���E��r��#��ڵ��zl9�R̬YӅ�X'����lK7�x�i�k\�j�ߗ�.p���[�E�y���������i9��}�R��sT�'\HK?0L`-��CB�'�<񀄣�-e*�L����211Q�=߫��0b����Sc�[RJzv=̥�m[7��}�m�J�z�Ib���������S��3̶Bޔ�ry����7,��D`�7BL��-��X�s �f�%��\���^��~(\��+^�-��̞:���c��f�N�V�	<�/���2s��Ts�:��P��0H3m�5�2X��yg�yj`����g;P�ή�Hsm����+��v$NO�6l����߻g�̔���96:RoJ�n���=˶�d�����'��(j�˟1�� U#��j�N䑵�����2��b�-�9�p�q��A�RslWd��&&�Q�8�`-�{
��
y)�{<�/Č57٥�� jO1K�+.����p��?��ȃ��"E,����,��8s C�C�%Dש�,I�$�.�}��i�t��ͭJ�d�.P�	��
�%
0V�z��^&����gs�P�4��Ҥ��� V� �\�⺜99g�nS��V?�QkUǲAb3�g3�������sm�Pg��,9��(Vc�$�C��+�r��/�|^F ����n%E��7u�E�o�D+I��DV?P5L��ℚ�;���z?�U�����Xq\*>����*lLN.�.��rE�4:ݩ�%�}-���ؔV=w%4r�,��(��a���e,ɖ.�P-5+�	���l��>�USg�N�׭�m�S�t���\r놌m.��HRs?{l:�X*k09\�Wl�����Q>cb�a[�[���`�I�f���n�:��w����ds��I�X���Q�H�1Ŀ&�Ee�S�3<��"m+�@{;զc�p���x��\�	7����97�;�JxG�MeY�`踸�PSM
�y��#k��27;�t��V,NL�z��b,���s��cY�Y��E]�CƋ���+��$�kD׳��Êb%SEB/mP��/0��+��	����	��m�:0٬433��w�ij.3["�����z�5���8�|��x���]�����9��62�MCjom�����R��k��J��D�����m�^����2�f�k��#���khʂ�Xt�i���i�|#*IY��6�B�'��S�qq���埜XWN�0�؁�j�*����Yۋor=����PL���FW4.�H�N��k�a�LOO�t
u2ML
>�b�|l�0Wr"'7�C:q6!j6J�&�g�ӪbD�ea"0�X,��fȆ)��Io��˃'��D��m�,�Vq��u�+,*�`������K��wc�<��}�b�\�=&�k��p;k��tt�Mϕa��6v4Y�@|���7��P!��&�	��4Fcjj�w}�9�l<vlr�ރ��3I�sa9��2G����K^�� �kvvnv���3#ev�v�X��>~|4�� a�C��:�[���.�WR�b�h�L��0�c�v��6;::zzz�/����n�-@�����Ҫ�۷������[�\:��S�)�i�7eÇ`�������M��=��_����U1׮��ןw�9^�|�ȁ�]皫�#S�k�o|��<�c�]��������(���(U�"��?�?���j�������e9n�RI��t�,\ ���^�&���mmmk�􂕍���janp��^L������u�뮼�7�)cmw�����?�#5e�,�uͦ��H�Sd�Wo�5 Aؠ���ǚA�Jgv��=�5��*#ϧ<:�3�pW����
��ަh�ӄ�.�A�V,0^���s�}��W^��_��W��
@�W���������YT�*X�s��$y�0�/���Hqp?v�J���dF������{MO�֭�y�(1C����ّ��c��ѯY�tA�4��/��LaEG�Vʋ`�ǂx�N�ЫD�x�{��A$�HJ/x�F���O����W3k.�h��C�wO�g������%�с��2�,���,�
���rE�($��Ł1>>��e�2T�.x�Z�b�U�y�r�x9��D�B�8��B%-�(�j�RH�e`�):��d�2�JBт�RȚ�<7Wu]'F�����jiV��)I�4��F�G�L;6�U���P�F*-�"O��������CNe&^�Ws.�x��"IŖY�`	�*��m�|�TS������z��7n����e��Е���{v�c�0B�=3�%0��t������Mg+u&̇��\��;b&�р��'�J� �,ۍ��n�Υt&�D�KX0�OFbȥ�`�>
�JɆ1���3��f`'{zz1�ԁ���DlBr	�?�g� �Cy/�}�g���D���tr�`I��^{囮����\i��7�|�?�U�f�Mc[�	@"qټ*��+q'7ߕb��t�ēB�F��X�K�U%OH�:x�.U�Rd>�*����n�_������͛0A��a��:x�3661:2n��|09YQ��=�.�B4/΅{����Ka�=�JD�X���r���ݖm�-�v���<w�����o�I�@���L��Ź�.��-pk�~^t1/�R�{DaO�w��]�
���my=kڱs���6n�ꩧ�8<;;�5��帶l76_�_��k��b�ȝ}	w]��!�yrܼ*�֍�o?�;KW���\*S����N"AX�Q��]8��-��B���<����0�f�Z��f�]J�4t\�w�ؿ��`=V���)j�T|� 2���!�R)��U��R�����߰!�#,$,Wܷaꌐ3�!J��rBpG��j��k�B!cf��;�ڊ�5��v'x�RR� m���,w\�{Y*ds8�e�͚��2%��|BS_/�j��I'���D?d9$�%R� v��: ���@s�~|ϝT�Ƣ_�*��˶C@�0*�&������+s�r*���.5ɴ�c�iR�Dp����7�몮��޺C�cWwWϭV�Zj�,Y�%[��$�`C�@l�0�q�<�#��#$� ��Kx	��؀���Y֬����]�]�<ܪ[���T���K�?�EѴ��=g���:g��ɴ�b�Y�:;5:04�.|U���.�c�|U�,�|�f�	��WX�1w;ȧ��V,gL��f����������Si�^y���?�h%3"D����X2�P�a�cCC��1146��rM+n5I����X��'@/�Do+#��W�hd��gN'�J9�R1��oi����"��@`�I{�L(N�[�U��=u~�UU$�S1*�l�ⴲ.Ԓ��S ��B&�q۶�����l��.�hX�mVn��
KdY����Qm*|#0�B����,vM�H �X�SEuǮ[6\s��pG樽ۈ�Mf�>甃wv�N\���b�9�n��P(�{t�\|�2"Og3�����F�&�Vy~�*o�Bƿy��� Y.�� �WYMrn�'R���N�����-fC���e��t�Z7¨��!��T1Y-/(Rِ#Bb`bS�	V3���S/���?�Yn����LLgO��B�=�y�w��ݹs����=}�g~2<>F��M�Wq�B����������gy��9-\��$���"tW����[��6�hkMm�׵�4��Y�rE���t{\l_�*�`<������u>������çN�9���*B0\c'�
IRRv�[t%�:�*ޥi兴=DN����R���,˗u���d`���*������2�(�K���%�PR0��H"�Hai�$ķD�:o%1��2k�'��,�i���J�������������z�be��0��ݫǧ��pI�<c7�&�[m_"�.����`E\AW��Un��j��"6nټm�6�S�XL,��ĺ=�fgf���cgϜ<�J!xcIV)��\>c�խ���<~,^l�6��f���������ոk�Ҷ��]>_��$���Ø�?~b"�͕)�R�*l��?PE�P�m`,�Pc1�
�MQ�+ ��Ʊlٲ��׮\�r�������n-�}}}}}�t60|�׎;����^dx6!��b� ��}c�Rᄋ����@�F��B+*�):R��{��֭���zzz`�v����(3Ci����(�.���CS3|%ϔK�dPt���%ӱy��7�x-��Z8`��%�Y,�8�C�+D�BQ�������Dn��֏<�h���f�5O��B�Y����0f��f���pk�Kp��	��`!嬪�E�BY[P_�Q@��6�f���zE�k15��H�bM�ƍ��v��� -���R&.4==��{�С#<a���)j�t*��������R��_�=�3�1��b����O<z��w�������;�6����5�=��!Z��<��T�ꭵR�9\���T��C�@�Uވh�@��v^�	q!�L455]wݎ_|����6VS:�mt��Z1K� ��i�����À������~4w�0� �k�	Z��ND�Ϣ�r4�(�H'��J:?�R�z�Ϲ����>���fL��Ww�o�Cx Q@������qz��0�Q@�G��['��^���~�
4����T&m��"��1~�y\��-@�X !���_]vCk�-��R����|������)��+o�rY��+YQ�b�'&��Z��P�P���B�t����u&�"Þ)��R�,�Jŕ�g-6'�:��566�ȿ��tp�f�s޷�C�Ž1Ւ�j`ڸ�k:��s�c���y��W^+�j��߸�������Q�(�&ZbYګ.Q��I(��D��>uN��Dђ���T:FD(1_�Uh_�6)م��"�B�9���74����O�9�le��[��Dx*�M�T�-y��I�X.-][!��Un��wuu56�Z̶<F�����|�\0��N�ٔ��y�eO���\qA+��P$���ad.w-�D,ҟi�66n�J�tv(���w���֯T������B�rX�������*�n(���x����NW+zϝ��jͽA�̘WUu54x$U&��!�f�*1.��Q�ck��Z�*)��ϥ�H�"ҁ�,��sH}EsZ�'���\(�HYџ��e�2���MR����h+Domcu'�R�Z�%�����ꞞZ]��|���o�`��.)I����Ku#d�f#S��[f]_0yK%Rd��"kn�uŪ��W]�����g1+�3O�3Y��P,�)��	���M��E�A�P�zE(�`Fe�� ��7����"��1���[�H��A��eCג����d����}�� �l��ڛ�Y�i���e��3�̅���@��<HUY5���CDZRT�	*�5��%�#_�����L�������<f&��vcX_p� AZ��v]�}v���Hn��N����ُ�y�����&ˠ@�T,U�<^+E{����h�� ��b�����z?�w-�@�C(�r��M�y���f�y�xK4�;{�������ipCJ�)K��0��(2�f|�C^�AIĔ�#����Q�j[[[W��j� l8J�X4�p9�6+�С���l2a��_L��/��'�~��!G6
�S�G�oڼ�j
���7�Hg���6䊂��"��b�m�.�Xr���W.�v���ݘ�e��@����s� a��'�z}�+�_?r|d4�0��X�X���O:�ͮ��u�W�f�Y�dL��(�Zӳ��6oX�q�Mrc����IgJDT�o6kyJ��W��у�`.%��\�y��v%;Y�1�"$�۪�Q1����-���`(�/���X�j���d޲�w�KfK�ڵ=�WӁ[Q���[�=�����̙3���I*�:��g,�#�ȭ�,��W�cZdVA�Q�.��J2.]ں~��{�=��uk:�:
yU�wV�ـ�f��O����������O�J������� .�8����J����̪"��m�SXu�L�:�F�Ֆ�Z���ս�~wKK���d`j����q13���0�ɤe�I\���?��-�\�dX���� [T*��fӚƮA&���ɋ�ھ�8���q�t,Y���D����Kb�����eͺ��ݱ��꫿{N�9�{v���D���[����X4�(�l!����DM�b��G��q�;::�t�m�fۭ��Z��T��P��0��6m���/������������(?,��W���!.�/Vx����"M�ꞝ�J��g����J#�ڗ��}���y(B�L4��<���a����<��ĩ������D�R��\���d.�q:�@u�h4B�����ȥmHtYfY����ʀ�-0��$�%��ѨY4���444�߸���iͪ�v\����$T����W}����?�G�F#�i�M�>�+�DN ޞ1+��;?����HJx3��VK:�-j��K�֮۸qs}]S.[Dp������z|5p�mK;��f;<$�ǦM[�;944GfgCA���)⋽1B�E�h.UeʕJG����s���}���,&%_*9�6Z�݂��H�R2\}�շ�v�����j�~��_������~���t������n� Y�=��/UV�j%/��y-
�'��#�S�N��t�.�@�o`�d�ج�6E#!����zӹ<���jQ�|�V(%P�t"C��5�]����{��3�������J��� ~�D����%���NfR��o}b|rdxl֍��N0H�h�%y:�49�mX`yru�5���k��uK:��vA�%:�	J0[��x�⽈����q�,:hk(�D��\ �d6Q��
�+�e����&%�"��̣E����w1�Ϡs5<�ɷ'GGGM�]�j#+}����,+J���T:��;}ꌪR��j��)�)�]R��i{�'��'r1������x/>٤Z�w��"+v�,�b�X,�(�l6	�(
��v_ϝ�}��/9~���d�s�V���D2T�K��f��k�\6��r�<R��/���Z�VR,x]/�h4�k�A�1U.[Y�lNG<� ��ee��_��o���_`��m��)y�C:��l6�H�F����~˖-�n���{E�D�dP �`��փ f*YR�Og���N�<}�T/\��L�`��2kU&ʹb��L~��,Vl�/Z5 �/iܰqM}]��Q��J`&�u�zd6f��e�9�0*�o�[��l+��+��c����?�L��\����B�{:��l��i���K	����|h�J-����|��nPeC�u;3�}}�-��9r8�Q�%"�$zcc����
%�J�Ӿv��ko������}����jV�9��	�_,{�^�TP&��|>K�^�aݺ5���Ӄ���##þ�v�f�V*�V�$Y,V���{Y��-s�Do��g/��j<]p�M	U]��h���T6�_!�K�n�K��eg���]K���Z����ș�����Ƃ��7KŖ6���.�f��c���-`����G����ɩ9�*��o�.TwP����V�8�b��U���RT���v+���+�ضuk[��;�����E�F�¼�@�D�õ�Y�r��[v�������W/9r:ɹl�t!+�<D�8����V�q��b&�agA*]O���ٶ��U7�t��7����҂'%��e��a%���oQ]6���_r�u7��:���=�����^��r�d����|�-V_8���m�����f������m��w�u�݀AX/X�`J󢑠%ޥĢF��|)�΀Z�\��{���>��?��O�GG	�&:؝Q&��7UoV[!��f�|v$�EF\I��P�޶��[o����klh��b���B^�k��A�<��RS������7��f��_������w<�L�mV>|&0�r�yQ+�s[�[r�����l:�J$4P&|3��m׮]c�ͪ	�V5YZڛ鬌N� �孁o4����b�_?h{���ssaL��*K%�i��	�4=`��V�#�|���V7 ��]6���s�� T���w��Z��Z����ToJz1��¡|�i�����ݾ�7�صb��M�|��?z�W/�3��B\���˕�K�O���*e-Y,�eaŊ ?�n�n��pz�C/�%o��N���u	u�î0СP ��_��/~�{�86��I}6�F��*"2�XRy�=/�����s�1-��daIK��۶m�zۦ-U���K�T�֍Wo[�~C�y�[v�F���7���+�䲹
mUR���Y��F&/�/ǊI*�b�N}$/��-��L���2im&Cs��5[o�yӲe�,>��\Ũ�t#e�P������5$�d����G��/d�@���B��;��I��~R��(J�|�Bټy�S^�~���ܱs�MmmK����D&���o����Q�yE�ӓH����-�>O]G[���X2���<r�H��)Q-ʅ[x��F�z�621�w��'����k���y�*徦3� �u���p(���|��w�)w.�}�;v�@x�y ��֮]���}���,ȸ-�b��T6�0)�F.	F��n�zE�*MO�4U��jqr���p�]�t�R���QV����
�>�q���֭2��Tq�l�����܊�{�<<=0J�w���X$)+F��Q�fev$%I�2���l2�Y��N�\���#cS��sK�vJ�Z�C?��Z�q��w�~�_��*�d������X�@_�Qq8 ��g��(?&�+����<��#��<01>G}^բ�f��siG 87
�9}��W����L�)Ab��څjq���� E������k�n��?Mt,�sU�D2z�ȱr� +ԙ/���@�t!�)XlV�I"ݨ�^�S�[��)b�a:kjj�Wsl����}}z��v{�k��ڛ���'�����T �LCAxN��f�Y��?<0X�r|��(���C��;���t�*l
�N����2��Y�p�/Y������L|�������'&�?O����xA7W(�?�w���bY�?�/�@z�
6��a�7�wu�mۼa���V�=�ʜ:u�"�Xb���`w oX�e�$�ryI46�x���V�X~�ĉÇ_&2yYb�4�-.�Y�J�!.�iڍ;�{�ч �G�ǎ?�H���[�k��P������P��om\�jŪB>�wa ���u�L����ؾ�}�s�R�d6Y�&D��$e�|*��w_Wx�'Z80��w���ijl	������X$�r-�X<��x�39���"w��ZY�������V.�dS{���%������߼���/�|�_jI�U=��v�u�w�� ��֭K��.\`�T��S� �7҉��nǰ����Tc��������}E����^���������2�2�Tۀ��ѷv�,UO(����=ݷ���>|?�~"���Db���"�(A�hMd3�|��7�	H��/�R�D���m��1.Kھ���=�{b�Bo{��8I\5���tv��r��{>��.����r1)M�J�$��*��7w�e�ͼ�2�ںƇ{b����������tX�M\a�z.tq*�ŏI�me����cپ����{���=��z��ɪ5&����V� �@��f@��zW�ݴj��믿�[�������x2G��W�#��`H���2ϖ�焍�l�w���={��Y��"�E��� Tց�:���U�P��T2M	ueR��X�~ݪ���߰�����_|��R�bSUN;�6���	��0�����Ւ�R^ж-��<��m����xV�2k�B|�f7��H�M5��Y�O��Ʉ�������U+p=�=��s���\��E���c��=f�=x�	pg�+�OE���ٵ��G?��Lp. ��I�s�"�7==�ty��X�2?�m^Ҏ����{������{���dr6���l"AN�D4����7���T�N��l$ZEj�_�>�/8�֞��w�������յ��4e;g3 32	)H�U8;_���7�FL%J�4����;�w����������_�c)�ͦ#�
o�~�EV;;�q3
�/GKS�-���t��M[�s�r�D���T@VTHX���k+��m��������}�70��ɔ���I�\F��R�^sXb��K���z׮�wܶv�UX��^��&��)ịeY�\�&�P�gsK�k����ڷ� V"&>;���8���0.3>TmH��\�,_�`�Xd	�_�4���{�s۵�Xk�*��@��ʳK7[l6��N	˺�1�]˻֬Y35�w��/~���~�*.��~�> ^�u.T�|����z�	z�����{��ݷvvw��j+�X6�����.=5^�>?�YX�2^�($���(c�����&>-l�W�d�J�\d�� u����٧o���@0�,�
s����u� �2)�6�)OD(R��XgW�O<��{�ݻߵt�R�����}�����_H���i��tr9�����5���X���c�F|����k����t�
�Q��	���L$����{�K��)��i����~`&�x}5��ny��x/��� �wRݭ�������T��x<��Ձ˾�?�Lf1�N�Z!P��˺h[��m�ieʢ��0�@��X#JYӌ�De�cO����yQ����-O�|�! #iLE"�ə@(nj��lv�������'fB}���nGgg���?����N'O�]ؒy�0A���澞+d%��z�V,_i&GS�p�l?�^L�c$:�̳�Ȥ�e�n��	��5R]�0TTT����P3
P ��`��eL��c���q9Ke-��r�T��%�E%פ_W6T���a�he�Q���]f(k�W_y�����X��/H҈�e������,�|1g%����21O�a:J,��XEjd�ӚY�Q+I}5>@^X��d�*�^)]9��ri:8�է?���v��8��\�����c�W�\�dI'�,���Qa��"I�T�7`2;����ٯr��w�X��;?��@��\,��0����C�O�o�r"t��w}��_��T,��?459c��Nk|)����U1�x��-4�6ֲ��B)��U�M���r�v����7����_�
��t��5Dr[<���pt����<����ۛ�ȿ粁������\ΤL�ญ���fX)%�,�ZNd8?���T�($�`�f��p�����=o5�y��+��qM��������:߇>��c�~�y�����Ó�S��� O��)"R�#ՌQ�qܔ�_�k�0Z��x��c�#Ot9ܵů�D���EoI�ȟPY�$K��s����/}� (�\.�b<����\��዇�L1�q�46X�y�Ŕ��VD�t:MK��'�lll���}������'Bo�$!K2�Du`�&�t����_v8]�lf|t�nׁ�+b�P�F�	��v`DX���Fv��˖U�,�����/|���W/�ۯ}���1.�S�0���AF�ɩQ���eݳ��G>����Y��p(4>6c�:jj}@�g7��/�a�7��1�dN�êl���k�kI��'?yf|* ^!K�������eq����'�����
ŊP6��%E%�r��%�w�d���Ɣ�H�����`���/���5�4���W�����3Y<,���r~��A\	�$�@�JZ���Y�n��?z��߇W��I��f6��I���Jp3�I�1�ɀ-��S���/�v�I�7�qӦ����^�v�׿����)�ݜL�
�j�B�+��f��o���ݚLeZ��|��׬��q/�l�������B�����Ĝ�?ڱ��s�2��g��d�vLv�@��Ҿ��G�ꪫ������g�M&�
���p��%�U�d��T:��	1>���+���<���?��G�[�h��D�5�R��&�j�
o���s4��	�䢍FA��Ë��-?��cޚ�/}��L�g�Z�ߢ(h�+旝+��j<��l��֛v�ܱd�`%�d�JZ�b� �v��偁+�b��H$Uf�f�ٯZ������W�������cB�"���/�ď�/���� m�U���[o{W{k�`�d�B&G|�(�syI��*��@2�eR��@#�����[7o����~��LO(+����b��ՉT�+���,V�aK$�JW�Mg�kk����<�����:��T�,�L�VF%%���`_�f.���fj}>������/�پ������ַ��ay������v���!2������=��?�ȭ�ߦ�,��Eq��n�ը��@�d"�+�@�6'U>;-�t:�4 ������V.��K�����p3�8�yhh�������DJK�H��6�����8��9������Kϱ]�����~�h]��W�q�"��Tez�:��#)YL�(����[��P(#��V��b����ٳ��l.�I�=�{�}Oc]����s��-^���h8���\�d��Z~�m�/���������=�]>��l�fI�u}d�8�sv�kA���si���7ONO�Cщѱ��LN��r��w ��f����33�2���
��N�0�333&�\z�A����\�����?����&�ӟ��'IW��Y_�����qK�l6@	G3����nl�ͥ��N��Fc�W�f��p��9���C����-^�\,%X� ��+�t�T�MOM	�ܽ|u粕����[��3ϼH��:l�e�R�b%���K*\1�~/�R���ЊLt��`D���es���9��@~�����|�A.&>By9�j�C6P,��2�.{��$�J�;z*��2xA��Ԡ�Sra:)YQ����J4�PҊ��+�ri����]�'[��:>������.5t��2���p�K����_��=?�q�<���P$�������v�].��m�i7_�9�lhI5+�U Z�T�d�4�6/Y����1���"�l^�93¸H�L:V�zȐ�Ae��@��Ɯ�qIл��_����o(s��9p���T�l�'�i�p*��@b�X��D2U�9);��JF�JE�+�l������=�����޳�RqC�u�ZmF:ͨ,����c�`�
f���ӳr�r9���_y����D2�l�YK%A�M��&��㭱X��V��d�O������L�Z}c���މѠ�]��
:kJ{%� �L�����ݢ��}�}���a��w�~=84*+�D<��7X�U�u	��P��p95vgMSK����sLE@2I�+��\�=4|al$��b�؊Z�"�21\�B����R�Fa��L��&���'���g��R�&��X
x���^���Y� B`*���546]��*UQd��2R���J����+V.�\�?pvf2h2��D"��D���l���)˳R�1�զ$�X��l��G>���}T3�N�F��v�q�����33Ӣd����1��Xh'^�g�99Q6A��Ky�bZ�ٵi���^f1*̍�%�WŰ^C�x�o�R�+�/Q6�
��/��j��駟x��z�``]`�bN�����d��,�M��E���*�P6�����јJf�M-7�W:~�0�0�?��UL��0H��9�
�*��?ú�����٧>���?�ty�v
 Y���K:L��+`��t�l�Ah��s����`vb�$L�SS��$����k���v��	�۞N��e��y�O�u�p���I���+�$u�����_����_Àh��bguDb�H1Q6}����f�`�9��+F�F}Wy�@�hR6��v͵��}����9`;�V������2/U"%K�uu^�;�$q�ՒNg������О�{zzp�Cc�DV5[�"��`����L �kK�2�T��6�y��狠(y����mI��X_���J�v��)L7�a��;�`�L�E$�M�%2�+X���$i�H��&��m��W��'�p�=Ա̈y�UҤ�����hǽ\BRѸS�_��	�J�|u����8���ꕫϟ�p��i�#�hT�]����;ͱIdy���&I$A~����~~Ǯ��-�����J�n�>Rs�2��B	�"x��%���<�I�0���m_��u�ܹ��)�M$I�BQ�_>�'����?�R(�d>������.>��w?��G��}g��Mױ�f�D8�|^�ƀ���<_�Ȟ,���s����k��##c̀�H$�p��)��H���6_�j��a�N��n���tN*�,d��N�iσ�������ɤUe"٬�u����ҙL,������=z\N�
}��g�ڵ---ǎEF�u2L��Ȼ�I�␗��nK�_׈�V�-�1oۮ��ɏ?^��&�"�mѱ�l!�h�I��NO 0�W*��ڣ����D��I�4�̤R���L��`cR������X9*%��|T\/L�K�jV��u0Q%��������5:�:u��/�499ɖ���c����b��D�K�o����*$nd�f1�$#�`�&وx}͵��E��d`���z�b��fy�ڞO=����Tpz�,��|.���V���T6$��h,1�QL�e+�k�B<R<y�ԅs��
�$����ճ���\a���DC�k��U-�-��M�t�����zj����$�����a�8�8��J%b��ccc�C��mm��z���d�ȡï��j<�zp����f��2�5�\WW��C�Ο?��_�rA�uŐ��j��8H@�`L�ML����܈��|yrr
,hٲe0��T�?�^�ED�B's��h-�x<&��h,�f��U+׺�.E��կ�u(��w(V���{�b'J�%Mx�2O�(�G����)]���
�K���g)�S��7�+N*��C����R���/�y��UC��AVv���WW[�� DH�9_,�Ya�,�K������K�6����zd���1qfz:�͊�"!���uq^̎]5'B�`���w�v����SO544g'N�x��_���cĆ�F��a\[()Ѯ�S5�m{����vS�j{J�>���"�������D26<>����bǥƒ�ʢ<��Ȗ^a�E��
B�2��H��M.�{zzj���g��&�	�d%�l��P4�M��qJ�k_������I�x?x�p����n�{��ׂ�Q�Y-^9o�f2�l+8�b6d�G��2�L_��s����&g���fI���?7�!���`,�oϊ���z�����j�j;��E"с�AZ���yߋ��Ԃ5U}�c���g���ɤ���@p�Б��m-"rg��S�N�3饝��V�äʼ�e.��98T�K��{��LÃ}33Jt4� ���Ƣ��0ߨ���[�5�)F���@?�٧�ɔ��L$f�%��?��̹�{�NNN�b	\�����uP���"k.D�:i�RU4qE�I�4�á�!#hɔUN;�"�"�x�^j�$V�?�x��G}����{f�ɨ�C�p8v�ȱ�'ON��5�
h3KYj�2���1�t��N��Q�s"s:�]]��'O�yPt���(�`�4�i$��L ��d�H��駟~����2�Q��%Fibb2��e��s#��sss������ѱ`_}�.`���+W���.qf��:;;����;Ȕ�d����3D
���cJ�mjnĻ�Bs�Hp���O}�ݻ1D���
��DN�dIe�q�333���X��������^bN��ӆ1,�t\��Ç
�"O�)�?���B �������|��K�?��O�u�6������l���f��8�����
�F�i�
���rd�B4�F��h>��&�VX�c��աP����>���K�|������b1Su_6C%G!|>�~�7�tS������,����n�D����*,�>Yw�耋�����W�[-VZ�:::v��A���;h|����ˋB,��iS�� D�(����!�Y�ٙI&A8'�j6�����G$��=��Q�5��Q���b��E���6�DP��f��&&'��G%E��GO���@� iV"���ߥ��bz�C���C}��o-+*�<�˓�L��e}�u��&Egj"�Y����6������ q�TjA��� ��*0_.�3�-J���Oe
�M��?��C��]㭯-W0M&E������X�ìB�b�� 	՜��w������s�pH'�j�	Sw��+W655���NMM!:�l#d��Jv� ���`<��T2��+4
�%m�w�~���4�I�R0�d
��Ҥ(�x|||:�a$��4��>d��^?c�X8�C@8v{�&��Rڈ�6;f��fz^Dg��Ә�V5�T�/��}�mW_����o���Lı��X��c���\
���c@1�Kh���7�4�	�0U��ph�"�0�����q�-�چ�������3�I�餠�mf���7�߰1ML�O�4���#�XC����?z�X$u����b�p����ё2I�k0���,<ښ�lي288��55���z�ǦW�{�	oY�UEx�� 8�X4��;���Y�c�۰���e"Z���>t�ĉ������u��w/]���!B.\ Z�`gU�T!'�B��������h1K�cc��P�������b��oF"�������	(0��f�bQ3��M��:���4!�@�c�3zI%%(�h
���?��߱�]-���1�,~2�3�Z�̓�\�d�2�+�V.���R]�<�����q��U.+��4�D�^�ɭ��}�c�~�#�ZM�����Ғ�F�����5�� T����Y�2;�52�	�����]�6�ꦦz�U����9.@"�u��p�SqA�F�m�9d��6lx�G֮]�E8=5��0==���C����$ޝL%�G���,V+�/����l�����y�22K�APTT�����j\�����b��pi ���<2�g�	�jH���3 D��~��]_�����	��R6�AD� �29`n��b��(U7(`�Kw-Ҟ��P����{Ϝ��s۽�촂� ��=>�䓟�Z>t���đq�98&��l�lhט0�ʇ��t��k{A`�ӣ�4�<�����n5�Ν;�)t�A�3���ߛ�<#O���;���/�ݎÇ��)���c������a�5��W��(Q&��F����U��t*e��y��x"���˓��ɓ�r���Ȭ(k�"02�{)�����?񲫯���/�iwOO���K�&�lp��g����o���d2��o^<�, ����UQ>,�����L�_��d����?x`?��H#l��&i\��mX s�7�i�����}�_m���@����s}�O�z��_�9s�ns��p�'��g�p�fÃ�C�hf2Y�z�`(kN2�]�ёᡁ!ک��������e^��+�5��Z�������Smm�媄.RGb ��g�@`rj:&�#�>�W3999�j	�镎���G �e �����0���7����/d�S�tWt��]O�	���;o��K��K��fX-K:���(c�ÿ�s�V;����ǎ����D<r������|u�yc�a�(�����pG�p|�v��5�"�<�sɒ%������A���>���<�����Q#E�*%LfK2�
�Ύ����ɒ	<&�kŒ�e����!�b�8>-�x�`A�B��r�[�6	d�9'mJ�"vMY�LiG���w4hԍM X���۟�����
���;v�-LϤ3�Dbf& ��!2F:�Lbu�p���5��X2�t��'���� &?80@y��D\�|%zU��a;"�%�Ȝ`ŤH���3�Z�͎}p�V||.�O����r�Z,���40n 0�P���3�����7��8�\�X`M Kڗ�������Y�|x 0�!c�3�ٙ
�]�m�͟��Z�F0J\瘩�R_���bw�c�Q�oJ��gϞ����.��p
̅�������uc.���%�g(,��9���K��I��bx���=��?�a׍�--f����B9_��>�LT�B/��GG��{u��}}}'����F��UY�b�D(<�f���p�@%�y��V�*��t��	�R2Yj�kw���"�Ӧlش��Q�6*�)�$Q�x<`�SSЏp8�(P*��3���f�� EX�XJ�d���x�5��C�U��x۶�\��Ǚ93V�C��(�֭[���'7nZ��������Ը�.� �|ll�B_�L �ZN��/vI�B�n'���%@��h��"M�l&���b�2�X<�HbmM#����)�_�V�,Y�fUcsKSkksSK����ڼ~���ΥSӳ���=wt����ܹ�P���2Nh�d���M�rq�M7bi>||r<����YU���0pp78$��:�o7Z�����DQ�b��͆�0k+z��ҳ�^0	6r�ܹ}{��h0W�,��X���{/���S#d�:�����q|&�0�?pժf��b�XLƥ�Mk�,9z�/��X���IZ�jթS��=JZ�f�G�K����R���\�R!_VMb.���h�R��Ţ�-���zjTKax��/��"�oN��\�}�����!_T�{�R�+,TQ������PU�|��_�/�E����Y�����YJ��B��/"�L`�:�Ɠ�����aD;������"Q����d���
X	4Y~�V$�ju{dݼ~���o�94>ua$(l(k�ݻ"���^͵���.T� ?�7v�����}�ȑP(�t:��W�Z}����07h��œ@���Z��,�o�8}ر;���
�T&���w�?�ߡL/�m��PIQ�De>uMxc~���������O����Z�x�0__OQjrbZ��	��E�G ��訯��{W����&ŞLFL���?������,\Ah�""4�#s�\��S������� �W@4>�F��G
N�w&����$�5<2����V�k����r�V��	lLc��,�ڵsdl���_E"�ɞ���b1�R�������oii��+�M�S�u5�S�'N�ΈF.+X�LM͸�V���ŏ>:7-ie�ݱz�
,/�ن�CHfl�TД�ʽ�ރ���{>�5�Mj�$��3�Uu��+p�K{��|}���G^�a]*%���h�˿|���ǌ$�e˖!��#�l.��k�
����po�tuc����J�y�M7+v]�M��r˻�9�O��=���p��	�-O��������=+�=���~6��ح�l1�{����0��3g1YԹ��!��`0���������9�����.��U֊v���Httu?��= 	g{,6w�P䕍�T�u��k`�uVv����|�ӟnjj*�K0C�q08w���'��VYې�����Ta^,�gg��!�<����e�}�~_#e��&|�e�����h�S;�ݒ��X�%�9#&؃����&��?��:�L���kEvNL׎e
M��pG �����V��7���Zq�G:|)�o�����'>x���{� ��Q���P� ��/��Qؼy�?�A�l)f)�,�T,��`���c��H�*%�$�N%H�^�`�N�/�7H{��9x3������747?�������̐xX+[��0��
��_��4�LJ6W�nm}衇N���Mŭ����(NO&�1K�������"�����ہ��|����1��M����?�|__�k�puf�<��!��^�,��*1�O=�Tgw�̗4��t�X�Wb>�l��Y��ߩ��T:�o��\j�B��������0����@��n������g?���r��'���kH@{
�$S�a��s�����]]�VN��1����3`}���A�B1�e)�]�A�O�>��u{��{V.��zeń���zq0�O?�4.��r�t��T�%�V:���Kxe�P�Y�QU�����ӟ��w���$ATL�X4
�ʪ���o6�ŒO%18��`��+�Q���\�D
�ʟ�	"����d0�}�C�?��?�	��Ȏ�t�<z&a ��]¬P3V*$6��z�����^��l������u��\�(.�X�<�Lvk ߅a�\�L&��$��gR���Œ6OM�+�dm��5v�Y�ʄ�T�V�v��mÆ=+��ۅ�*�Xm�o~�������O�\~�����
�S+*��ai8���j��j��o�6<2��ؚ��*z��w�U�I��Z"+����NcvRh[�V6TN�<���G�����i�bhr"	���g3�v�r�r�5.$؏O��~��իW~��?;}���=��)T$zR32��w�^o�Ȼ`�g4f"��fs���u8
���'H�F��D����̪��]����='B���?�<���al�Fc�+�bm�Y^�I*�R&�������Ŋ%�n7���#��� ���X�C�h�#�?���W(&ַQ��$S��%�X9@Ɗb۾}��.����~����K��,�77_���9T*����\�������g\�y�bnulv;@0��'?���-[��@��wy܀Dg����G?�=w�>����M�Y�J��lRmv��Fh�)� v��d�:(�Y�XT���b��`<�2�2�m�����w���l�7�޺u�-[�Q���a*��7�q�����~�UfS��F�|n6�F�jU�������*#vPwd�Pd�k����������E�5p�,�H�U���ɩ�f� =Òv{�X�}��s��9��`�1��o��U �xO���N���>Z_8d5RYTJT8aA�L��l������҇Y1%R���Ƨ?�����ry Q@��m�&Si� �jw��HƓ&���W�r����e��	V��X�ز��R��e[��ett�̙~�&�Vb�q�V��W���}��?$199�t�R�����7����d��P(�#�c��QP��KZE��.3���F[ԒD5$�����I�A�1��B���o��zϜʁ5�eeA��#�Fn�L_{���i�ZKE�d�gS��ə���������|�27�XL�,�r�����#sa�W�ٞ�(�-6�H=(ˀ_L<���IZ���r2@��ZQQ�_\Z���X�����S�������8TU}�gff�3�����ɤ��@Xp�>vRK�����:�b��g�s���֚�%�;��X�6�""bE���<�)����=����#�R@J�g�D�cǎ�>0�@0�b*q��V������/%�QN?K��J�Z�b�)�U�!E��ٳ��_�%R�}&Ь�`���v8����4i��;����Od3�ق�Z��`,��p�@������ӧ�s���\pbr���Յ+YfŘ��G3���?��r��믿�p(�uA�L��&��g`���={��~��G���Vl��I�t=�΅���S3�c� b�3���Bs�T3�Y�o�Iҝ.8\O�ߏE���#�D>H�7E��� ��2�	��Pu����~�P�����Q�848t��q����b��l,�E��?S���i,��7�ve�Q3x���>����L�X\���C�j!�LY.i`t������� &lȖ'���Ӏ���a��N�9�f0 }�.�??480;H�R����f3�.�]�`�|8;��Ra��RlU"��lY�S��Ԏv wI���io�����x>�Dg�ip�`pp`��L�S��ra��T*KY��\>�xc+��H�+\ơC�(O��<�f����h�[6g6� �A�Z��}�={>�G�G�
�$��YR�R!OM�"Φ���lhltrb��4	p�FJH%Lܚ�ns:�0 n\6�円�8y�����a��ʈe��v:�k�����V��������sǶ�[j|�M-�6�C����ţ��.�"!���!�F��r�7����$0�XJ�-/��m�e��}X�c�2/{��!f��Maa��j��:�������ʐ`�om�������mI(z<� CO�S�Q�����"
(�&��*+�TXK�zj�U:%6�3�ёс��  {�l6��y���Q��d�:�B鬪���[��f�^�d���Ra9�	��i�%̬a����%<.�/�r�}��{V�c?��/�[�����E�눕W���&o����D��_����V�w����vuw/SA,f����bA���`����Q���ڕN�0���w���C� G^x��GU��¥-4P�/��X-ֺ�&��Z�ҠH����.���(&QU)g88���Ԅ������"�"��1��9��f��N�8��+��n��ge���;��?���������]��bm�K�;/�4�����K?�?z�F��H"�����O>�d.�y�w/'S����������~�����.\�#l��6���$�L�
�����ˆ�`�#R��V��-kT�Y.���������gm&+�|r�Av��ƪ�D�Q�%�v�����\i�lr��P x���g��RH��慲���/2�4�_�֢�������I�0h�"2��,��7̸*��m4��O�Ler<�T4��}��u֗�WXU�::� �LMM��B2��}G�Y�
�|.G�z9�ʒ�n��U+W�dEA�fw��LE����b&/���'�g_�wP.�g�r�һ�s��{�xlt�ŗ^B ��z��K�h'�$<�L&(Y�"f�0,�:_-" �x��ef�	��A4PA�g��%�Qw��w�2��^B���6U�q|�����K;�=������t/�Ra"�d?c���I¨��"R�&94`iI�'<�Xջ�JP����M�H�С$�\� `�nI`I����zn46���+_i_�	��� `�����?�	�1ctDi�
�)�g�LOO���������C��[��v'�M�iT��kCZ��5>>�w�>̅�H,^�F���ɭ^��ӟ�L��!��N/�Xzf&p���c�^��;Q��"��x�-�y��� Zj����9�@+Vl�f��_�2'Ʉ�DInin&�>�G��B���{��!����K;;x��R_߅g�y�UU$"?�xf3)cEOaJb�b1�KV�a����>���VA�H�r�Ht�f����o2�,ϙ4PoPjJ��d�aQ�7��O�=�V���R �����fIVt �U�̙�_~���w||txx(��!��(m�>���|W�*
L&�ߵp4�ZԼ��k�J~�@
���b�`�"�BI�T,7���LK����n�u�|�S.����TK2���%��4&.��L�L�����b�cl1�@T�:�� a��� �'O���+����Q i~��K�AT�cX�z\qK[��ݑ�QnM��N\��ؿ?���ˤ�S!��L ��2��`�I�	�	���x�E0`��U����zt���9[��)ė5�D&@<�-�7=��O��۪&��<_=�均��Y��rLr}���V��D0��M�� � ��>@��l�z����bY�lى�ĳ<�PlͲ�,i/?���c�=����%*ڃ(��)���r�1/��ǁ�������L:�xO��pd�hb��6�׃����1�a�~��EjT��h;]vp�p4�!K���|�3�hnn��J���(D�m��f��ё�������g���C$��O%�%�iAÈa�����j�l����Lp+�����D:���ZO0U"u�J�O�@Y��0��Ɲ��}�vwM<��fe����6;~���t�>�J������(�@u��}X��Q㗩�qv��ದ�r�E5����0Sf��E���ԙ|��q�ꫮZc�YY�!�S��*�rĩ��F��FL2N�+��.&]�?�lS�0"v��L����F�9���9�a�U���q��M-vO4�I�8<^���*��h�(+��u劎`��f��sE0��Ȼ1VLE��2���|.�b��k׭Y�zrzj�ޗ��]7�9�,�JlQ�SR�x�f0j�B���'E���˻W�t�ɋTLA��f#g�^xm��f��r��8LV����c~{R�h�k^<t��
��\p�ı#��պ��h3CY��cfz������7�����������h� A�;�M+)�J�V��h*U��3N����������$���ɌɎ(Y��Hw�@ ����n��w�}����ν�M�"���f����o��{�9�����߹v�666������g���;�I˿��D�	�R��SU�ۣloo�,�����>��ř�|�;S�V`��軋J{3�7&l6��$�)���"wI���4��_���������Y����*���v�u����kg�x㍁����/|�������C��k�U���I��u�L��Ņ�۳l�����Y�@��	��ւ��{�}V��?<��g�<��{[�� �mބ������*�� aS�f��֖���^�a?�k�Z_۪k>�v�)���k+˄{���$�/��q6X'g8Wʹ�����]ZZ��?��e2E���Cb�y^��1K&�p|�4���v*�����TJ@�>��VWA9Xc�%$t�;����s�5���P�#r�������:"�*;�Ѹ��W�O�_�����<�8��S��|�b����2�B@Bwg 1��z��Q�U����0�a]��˰h���%5[�]p��>��#?0?��� Zb�a�ň<� &���Zͼysz}}�R����r*�2t�l��@k�zUV�FY+W������\&=y����_�2�b,�6�Ԡ���Y:=�g�yK��YY�����n�W��W0��?���}��T��A� �uΞ=4��XI��	׃��u�vM[ͥ3 ���S�R���{����[��&L�f�.j�������N<�H���ˎ/��z��M5^Nv��	0%S����b�t�Ƶ���>x�'��2L�P�a��q��tZ����R�X�C�����M����(7(�ͅ(��;������D�T��#��w`vHhax}�ѓ'O
LS�������3�\�|���:�q7LCq9��S) s��]c= �1F�#	PGY�;�x]��J�{�G�~��_��۰n�~��w�0���I�����?u�m5A�aڠ=�bt�Ӊ�p�����mzLc�܎tf�	�NEL���§z��<x������v�'�<!C700��y�& +�ұ�X3���#������>�?4����*,2j��byy9��{\^U�Ah˥B(�q�T��j�fuM��+��R[ۛ��X��?~�o>RZf�����o���۸5JVe����0x`����2����s�;v��uK�I�%QA<�G����]^�{csE����3���n�wj��ZÞ�5�1����b1�S��B(z�^y�[[�����`���t�R"5�Sy�� `m*¤}�m����$�ۙ�d�۩b��G�P�-w��7��"ۢSĚ��FǛ�YG���?�Q�Z���*���%`���-\?��):,C_��Tt�����*_S[0�*�N١:��U�1w{+�L=���2�U"g���Zp�
��Ԍ%c����S�"���$�ޠ����}�w�>�f�P�U>�+q�i�t3�z]�	v��c�>|��nO�4403V�O�ϊ��'��z^y���ťT:gW�.��-�@�n�䍛X]��x?
C�A �M�x����o�Q�!8-d�\(�/#�%7�������y�1J���^�ڤ�'C�c�+�*B��ʚ��@jX|�*�X� �q��b����Q�9 ������^�N%I��1��'�v#�h�Ȳ�B�D �c�)��2��R\�P�T㱤�*�����9�AY�Y��:�Y|���M�
 �ƴ�*+�k6X2j�%
�`,���u��g��6�{:ݡ����o��ݼ��P	̼��+.T��8���`"o0^i[���l�������}�F��?�'5=����旾�B8�<����d�7�xS���h����U8XQ�,��ܞnM�vuw(.�+J�;"�B,���'&&�=T�4E�W@w��O�f��$��?޹LU$R`��+�s7�_��nsy��n�$;�Յ����S���������W_}5�����-S �0X���a�b���v���������-��ƛ���?��˩��tӺQ�ImͻR����ޅ8��[�{�_w�Y�e�_˜���SO=���omn2"��C���3g�;�H�I�9�)�R��R1_��/ ��b��<��?��d��$sl$��O�Yq8�:�������5��[deA�3%]/�j5�
p�P̲�4�����$Jn���������dJ��,M��FN&�Y	EA��և6�v��~�!H�z%��ֳiw$��|��?�Qv�$�`ZW��U��~t1��x=�Mes"m�TQ��_��>�:�G��D����IR�"W���!�Ԕ-۠�2�/Y�5 ���m��u+Q����Vj{mcb;�Gp=kP�t���H"oӎx���!5t(ms���%I�u���p$�p+M�&��Kuj�)�f8iX�/:4~@�^A̽�� �!B#.��m��������V7��%��aZ&^��z�@ �+����u������C�b����X9�H�z ����p?��8ߵ�o�5��׾�5�gaa��}ǹ����,�<|E$D`��3v�η��8@$0\����Z�?x�Pow?�r�־�a5����K����ď��j��M��,��^�Τ(�v@0<��Umn����z�ʻ6�5�ህ��6��i��ӥb������C�^!<��"��,{L�Wk��%4%0����gϝ�-/�Q 5nJ�$D s_��!ݧRI�곳�o޼aR_aav�#�e����)���֎eY*�����OA����0m���j	?x���o�L�>���a��1,��qS��@?��K5�^-�
x��nTcyy�w�9w��d�+m�\[*�@x����ۛ<�䓸���N��U��@Y��9����g��t�Q��u�$��}��?��C�`6��!��I��L��kW�J�0b�{eeӁ�ru9ŀ�b|Z$�?���D��B�?�7::��ڊK�\�0�@�X�&NQ��1A��X����_�:X��뭗�nL��4-Ve';��F������gaqN��nO����$�@ɟ �5\;�n��i�9����,��F�/�����O�I&���%�3���v�c]����U�W�K�������w6,�԰��X$�g��I*0���r5G9�9Dp��C�l�L^^Z�'A\�(|�s���/~��9��"����^��#G0��-��℀	c�ao��1������u*�"�Q�J� TE��+��y-�ފ��uC�%	�Τ�8�����G?���&�����F�V��T:u`�}�TT�a�?� �ݠ�up|�$���˗�w0�w�+U���&�L*kh�mR�]7WKG;&wr�:���0S�?��O��	?��A
0���L�ۖY��w�����p�����x܍&(G�.�$AL�j�<��ֆm�m���0Z�4,�/������x����������%���7`YX��i���n�>����ٱ$��"��`�舻�*u:��%�U��+%b\�;�}a�׫�Z�kߤ���ʔ1H��4�$�F�E�|�@sD��TC��z}2�pjZ!���˟���%9�l�Q^��n_o߀U/����5JWƽ�q��ݐH������s��ч��%�Á{��3@2Ɏ��}����71V����G�ǎ��PwuOEY�M=��q��H�,B�+�o�b1<��#����˪���=�;??�Aa����x�n�Dho��p>J��T�n�F�����l���caOo8�V3Rm퉧�z�lعBv~q.�'DF��^����~���;���(�fɢpo�jQ��G����O�'��A��.��t�^��3g�`��x���^��/^y����?5\m��ӭh��4��;Ë��y�������n�"c��{�&��+Q/�!��S�%Q��"�F�v�R��?r��P7�����H�=}�*��$�a�gV��T�f�\��Hu�\�\n����C��Z���H�jX�+l6�hK�����K�YB�����,�[�6�*<t���V�������5Eg�Z�?9op�B__���C '��Non� G��~��G�O���Zx�u�p�C��Z��j��(�R,���HO8��IM�#Kdb�Ma�?��!�O�}ŚQרa�,��h����EA����%�����L��y�*B� ڢ`�rP�CQ��.��
9|'5�5:ooʶ`}:�U����Ε�IrBޑa�o��/�:;�Wזq�GzR�G�F�A��!�\�\�0����p�Mg�?�AGo�5~���jݺ0���vJZծ��1�G��<x��5�aɶ���0ۆm<x���X.���eUB~���<{��T*�4�I?ZU����P(�k�F���s�Wo�B��H���.�駟�F�{���pXX�[�,a�@�P,����S�Ac�}`��dKW_��@�s#��}�l!�:A.n�ذt������ޮ���J�������Cp��E?����J�j:]�?�y�e^' �:��q������ɏ�T]�����?�e� ����N�P�m��xqpp�t����7��~J������!��Z�6mo\�K��t�6+K�>�l�"� ��^�o��J�t6��栩+X>6�6�Db� �h�đ�F�j6�Z]�T�P����ɲ���45}�V����1���=]��TowO��@2��r^\&���k�ҍ��#�y\�A�Vw��t���߃Y�5�Z�sR�F�BC3[h?��g�����V3��r)£�MK׮]�2�0Cg����tc<�������{t�X���z�R�e����%����Y .����:�=��_�����g�+�S�r**�O=�\k{7<��F�/��,5�[�V/�WW�����`[<�ɦ,���9t�Ș���D<�ϟ>}�ƍI�r�T����΁#�uvu�vju���z������bu�*0?����u��i2/t�����1<qx�M�`ʄ\��ֻ�۳��W/�z����n��R�`�v��k�ЁÇ�:N��������T.�|n��s锡Uᣄ&�
|������9�:��-�7!�#e��}Ç��:*���q���:Ґ"���^�Պe��ݞL���1���|"��n�20���UfR\������c�z�>ARX30���pϩ;�n�;�`c��x8p��G��n��l�MS1p:�7(-��-R��fVQ�dm`�W�F�T*F½�D�����Ֆ��7�����<c����|[K��­
NA����~��;��) �Z����Ӓ�5�Z-kd��z[K���q��Q7�FYL�m=5�B6�S������:.F ��/ry]�Hg[��5	���t�������R��H0��{�g?�c�G{��,Le��nӪ��`k��Ζ����s�<�G�n�[	�JY&UU��RCR����	���v�M�^�^��se�+$k������������|�[�L�x��W�6׾��/}���BtԒ��ݞ���k�%2.���Y'V�E-��,AAٿ�رc0��K"y2;E-��d�y00гo���9ةl���J4ٱ�^�g�MV}Cݖ��1��y2�ٰ� �j(p��o}��w=�:�G��-7�d<�!��`(���2q��YkZ��*��-��!ǐ�n;�M���2�����cltp���=��ސ�������_a�����9o��̠����������T��0SR�9�hyei�X�!2�LN�S�N�:(�35C�C{[W3����\�-K`OQy����'���`��R�1"t�e5�͏�H��'���ve"i��4Qt'�]��)��￟�dq?�`(P˥\6������g�{���c�{*5�ȓ2'��Z�p�;��>�1�t���U�'���~T~�5�p��D� #��K/MNN~��_'TI�|�ÿ������g�I�d�����v�f����Zfg&�\������݇�v�d@�ގ���V��?\��%.j�0k�6��v��ZZ���
P��'�F��rW+e�4�A�*�MŊ>�X�4?�w?e�(J$V$9��J���#��v�&�±��^��֖ĉ'��f�穻�-��ι�W�)*	7�)[��l:�Bm4z��o&)$�1�S1���Ae^{.���|ʮ�P�\���{�E�п�ի.�˴��Ǐ���bM80��'�M���������5�d�����G�T��$�gwy7yjU��i�v�mX��-ڰ����Ol�u�w���@2zG[' ,&�5�1o޼~���������l&��ڂۜ�vKTӰ_y�����a�-̻��dWb,��F�v���T�d�v\%������rN�܋|\&�;���N�5�Bҫ��
���~l�Z�zܮ/|�s��0s�3�ln�R�yM�ʕ�j�A��kk�QLϸ�v��Ĝ�V��m��0�������;�J��h.ckc@˕t`�e ��Ο�ڤ��_�2��o�:00ВH����?8GϞy?�����nߞ;s�������8X��7?��w0�dq�rC����^�X�L�:jGG..k߾}z�>s{����r�v2�CA�ǡb":1ep�x<��d������� ~E�I�XQ�d2��i�D!�t���A��n�~%�T)UE�7�	��\�_�\��{��q/o=v��!X.�w(�?��.�/�I�������Қ��|��sW�z��w��"ʬ�⻿XixO4���9:�$U	,6�Lh��`dtZ�1��~\���P$��,�<y��ϟ�Pw�6�W��(s�m`���s�jVg�õw̋2�f����R�3P��6�jq/��7'nޞ�,r�H(����?������3�@<�Ё����߯N\È��R�j>��{ñ8�Ɔ%CX�n;rt��6L��Ģs��`�$�x*�"��z��8�ꕍ��K�>4k���}������8~���m��aX�O����iY^��=�\7Oi��6�2�����K�L��BJ"u�C#�@$@q%�c�aPP��c�dYL�G��"��c-��vj�|��������n����Z������z4��Ûw�aH�>w�p�{"��@�)`:v*�d�lؚf�64)�Pa�j���y�(�PQ��
��ɓ�p甦<0����.^�����k[��jS�E�,p7� z�}�F{{z@�,j\F&�Qɤ�C}������h�[�� 6%'���$_NR1��޹��=���ź���������X"J�~�^�f������l#�l4~�#�ȦӋs��������y�|6�,���Y��i�#X+\&���}��$׉��xI�u�:���.,���ˤ#���8�F2���޾���~����W7��9}����2����p��{��O޸~��ApW�E��;;���7|>=�Z�)Q�W���0>#RTkV��'��Z������LCt�:+��
Kg�F"ϻ���uv��W��֤�H�����4,S �mڽ�q��o���&M��!ڢ�D?{��OMM��є�I�W?l �z��?8?����u�D�-'�;�>��o�	�o�-锃�d�����w���6?}+�^U��Ox,gE�;q�j\%Y7*X��Q�t�<+�=s�VZ<rdAgGNEv���&t��u�5j�jRP���-܊�l���!B{m�>��J;M-acy����X2������G�7�:��!��)V��IWqhh��-�������������G��V� ���b���5��D��8�Vg�����O��mQ����5�c�l&������g?{��	��k?��~��_4Yu)�ů�Ccո�������`�F����/��D�%+�e�(������2k�8�����r��K�\_YYs:��Dls{.���*�֍��P�x<��S%E�����<�a��
-����daf�S+��/��'�V����-�"FB���Ex��}������-K�b�������V��["C�}�r��R��������X��3\	~���e�yVɀ5�t��y��� L�v8c���{45ݢ]�&@����ζvИ�{������s[[���NcP���)�=�QӉn�6pKc����R�P �r�d�JL�{I��#N���
e�H8X)ө�r)W�*�`?��3�������M��vaee����Ϧ����ͪV��J��8���4��$��%�(o�7��"\��7HƊ�5y�ӽ,I�� !D�b)Oɐ���p4��E{{��~�w��������������R��l��f��R`��[[�Uh�'��,��\(�ԗڏw�_]��G�_�dսm�<��W(�<_]���J��=v�_| r���/������яf�n���O}��@8�5�v���G�?���+L0/�|?��ڊ� �ԪRsg���A�9�4�5� "��M��� � ���U,�j=���Ç�KM��Itv��a��F㥗~���ם���+ޕ
E^��ĺ�5y�#\[(���%�S�sg-�á�J�f�\č�" f�A�5i__'�Y����[�N=�PT@ɕť�Tnqy	K�ܩ������ZZX 8l�:V@�I:������ML\㠄q!�����IW	�h$��Ts_� ! �L����&,Thzݰ����k�E�q9�o����/��M��=}Z�͵���� 橰�N����aB�S�G~=��*L���;:ں�:��d�6-�ٕA��n��h+���+��񑧟�Ky�pͰז��G����{f^�k�`�F����L^�6���Є�kJm1�.�����>��S�X�̖ �$Ut(����Um�o˅x"�?��ر@(Hz��czv٘�}��;;[�}������Z��Z��L�1ˤ �k@)Ar�D���En*��aƣ��$U5t���
�Jc�$�6��B,��+n���F0�S�c��U�*.�_(f$E?x���kaiym}c{+u���^GGKCl��R�N��`qKܚ>��Bh⒎=:22���JME��b���:�V\����+��醈�G��C����� ��/���Ȋ㥗^Z]1,C_Z�������#G)E�t�W&&��eFSa���[`}Z�h4�?���:X~iGR�:����q3�����r��u�<���b�'{��������H$ZF�{z{�_�.�w������&��HKP�D���cLS,iik����)Aƪj�R���X���0g��B�X.U�.o]7�����P⏉������������L�V��-�ᒎ?��b-�]�D��->2:�ЩG���o������`���B][Y��}n��-قK�����]`���3�E
~�ήG8Lq�\)b�\�z���_���W�z��1���lQ�k%�Թ�$l$@	�$h����-sh꤄Bڕ��˼?/B/qy����Uӌ�u�NզmT�����q����z�4�(%/������R�zz�/����������������O�[.�/���k'�?�liC�RT���	�5�FK��\H���G�b�};��ΪX�^� � �ڞ��U*���ֶfn��;:���B�cM �T
�w�⇗oܸ���$y��qg3=>�h�4}��z|
���I��e�X�8��n����k�/��F��#QSz�����V���d
�������h���#h��Ι����O?=6>��F��1A�ݖ�XU�z(ĸ�N�_�;�?�J��D�%V6W+W�A�F�����E��~�Q�7��_|�W^����U�\Dho[�o���?�e�Y�oH^��+��7��������t$���@�X_]/䊘��_���y���YX\-I�����R�x�- �ܸ~A�@�Z�J�Ѻ���rW#m֜���[��X4�ln}jrm��F��B1��FX��*k>��?40x��Lv{eu�R����n�&�,��F�'^*,n�����Z���?�������6e}m�H�mIb�2A�>�����;*�.s���0(��������ǎ��>�6;�:�\�V�`L=��� �lmo�}��Tzk򚄁5�ME;�\^��n�����x�Eұ|���A�	��%�f��76֋��P&�Y)k�D��%A�*k+˛����3���� �`��=�Vc�:h�s�_@��*����Wx�� az�7�N�hڱ3i�GV�9�m,/.\ ��<S���(�@2�
Ȉ_��{{�g�|�@[[�Չ�l*��`(0�������)ds��Ɏ���i�E���"�Ľ���4@1�+++�t����뀕�r�����s��z{;Ñ���Rw7e}�{߻u�>x��eL�[��2hQ̤RS��7�_G`������M��wE��VIE�#2Ϗ�!�����m0�`�i�w��p��ۿ����w�c&[8|��O}�xey5���^|�g��{�x�./�C�|�mҡ�W4B���&Y�w�N�`)������@,A��x.~��ʕ+7�]'uf[���}�'�W_��O.\� �/K.���ґ#G0�7oބa�������\��hfR�x$�� 6�/�8��������Et&������K���eT,�y�ą�cp6%��k`Ž==�?�@��ӧ�h����r�t�4.�s��^��ݞ��|�\, �b��)u�ɏ�x�n5IͦI�xT����l�EÅ|X�!��׭*X~,��"����l6>s�����������_\�B}}}�x�V!�,x��:���XK.�vttqe�=j0i,��7pN�8�~���t^�v�]M�sS��ҤR�TpG�;u�T:��I�[�����o|��m-.����Y�l:T���q�h��7���~Չ%
b����w�������q$`~��surn}@B�|�(�2h+�������/K����lN���)2��������&���κVZZ��j*��@Ψ7��b##�j@�+R&�D�y*X��z�2)ȉ;m�qaz����\*W���V��jkO��+W����~���vc}cޥ��mnzr{s3a�adQh�A؂�G�+�(�A-��~ o�{��ddWj���T�4M��O�aq�e,o�py�[��
u&u��X�,ͥoLN��6(��F�������}����k7�ORA�C�dPE�������p8H)M[ޅR$0��S���8�����f$%cV�V�0խ:[�q���U�k�ix�l*��x��C����l��Υ��a��v|���������~jj����}�C��T6��f�{^�."�,..7��N���d݁���Zs~~�?����������WI!���*��.�L��������ҥ+��=��w"�݋�2E����?�7����V��@FС�d�������㘬��5����bT�N^��V6R���s��1x���������̙w�]��rzO�pI��W}2�����G�ƿą����u�ɧ�&�ݰYc�&#��V�ߞ_�e�>w��[p��P���c==}� ���\�
KHe�W؃��������b��.���~cD�,�?�@v�I���T�����pO^����[Z�����#-���4�������rSu�
�������8?���*����<����Ǳ���h����Ň�G�9�`��K��Q[��S���s�!�������	t{���w�}������ �}��ߞ��fGw`\� _ð�F��������G��_����R��6��2;����b�d�UuH�@xuuKf����2xF>��";=n8orr�%S%��M�.�{=^YXE��=&($�#4�O&jީWa�5�j_'�x�HՊ*�r``J�I���&��jf��q:������e��킉2*���ţ�b������mj���p����S/�o���o����� ?�l����u:M�0�<��C}}= y�K�pC޵�%����I@X KؠoÒ�C�6 )��z,�=	�=�6�x��ek�z�,J6��V����O�����#�<&����ގ��S'���=w���ި�4 ��R���!ol�����6% ,��|�LP̩:hgݡ�q:��mG�5ր��HPU'f��I;� ZP�<|�F�)fo�!����k�&'&���н�@ ���|(
/.--e2@^\S��Ӏ(2�3U��X*���������N�HSضpI "��T��:����.��v��E���Ξ{�7�����g���?��_��2ee��+�ix/��˗1>---�3��(�6���� �ůg/;��}�>ņ%�����[C@���1�l�r����a�ӳK`_��{
�j(�-ٶD,|g�\ø��^�ra:�O�2*�<f�-0�ɋS�8�u-�9��c�p��xnP�"Xh<�y�q��fcp���3�����?=��o��}>����Ԫ��\H��yRU�Ȣnhx���p��^r^ƻIp�C\'6��&`�X	XE�b ��� �c��u��({=�/�˳��X9�ɸx�&j\���Oby�O�&Kg\�*����<Se����z�V��+T�M�d��o���W ��j�ݮ ȡe�Nw kEpŏ�ut�3�k�+ހ�Z���(Y�BO�O"����w[�B]V.6YŠݪ��C(�L<��q��l���x���n
d#_����%�iӹ��с��+���J6��Y���/�$������ ��X�~���m�P�@ �:�;����q[�r�j�]�R[�BN��\�]�mj����jes+u��՞�ζ��Kuh��$�UI̤�n\o4�d�t͕�'�m�F�2�N�ʕx�~\ I@�� + �L�o7�UcV,����:k�����L&���G|O[G���ƙ3g��G��w�8�͍m0�g�y6��~���� ���`jL�5�W����$>U(�yB
�f F���r9¡��4�����0�$��v��,�;�l��������0�x��a��kW�֖6{:�^5T+i���<^JO�6V������r��g�',�vX$��$�5zEU�uyӔ)U�S'�ZM��,[��L���$���@=r����b�\�TG��+�ҕ�ʗ����Րr�����>���G|���Zj�֌[u8p�/P��`%�REtЎ3�Ҫƺ�,Ϩ������:E���,��p�%���j��tM5
K����\Q+E2�^�̝d��3�v͟K��HDQ�����#U�?"4�RA+�
��N�@�Hz���������(�K�p �/YM�G���w��o���W߂MŒ-��N�挻�?줚/�%-;1�Λ���5���n�#;�ۢ m���WLCJF;&�\�r�r"�������a��q �c~뚹�����?�v}��#��O�>=k�,����$"���Wޫ��"�;�D���,}r�a�k##�Xߣ���pW��I1�Qka=3?;�	��~��Ȉ$X��7_{��K ��z!�mU~t$����,�Ĥݭ��M;��V��7�r�*=�˅k\^ZO�q������y2�f����?��>8O�����w��������8r��ɓ'�R^����Lom�����Y���n��衃�&'o��Ņe5?��t� N&��N��t$����g�qE�[�J�*�R��ޘ�i�B���پ��I����/��R�@����dS�p�~*�h����5����z�4V�U�zE;
�i�� �ng�[��X�j��5]05D�h�Α�$�s��}vѢ������T. �D��������\.ۦn}�]�O���r> 8:���'u�.�4�tp=07�pU~?�Tp�iD)bB�"�k;ض��� CÍ�o�Z�'�$F�����W��oܘ�~���c'c� /�
o��׮^�2==�_�,���d,����1���LUj�MjˤЙC �傘����)J͠�ήv*�g�AG.�Ύ���m�{�XJ�2�o�=��3�ꚑI���<�?E'&nܼy�HD�}��a�`j�H4�(n�I�u\*� 0�z�t�D|c˛�0�}����������gϞ{�'�����U�ɣ�?�[_����?�˿�h����E��F���z�J:ѲH
�L�������(���i����%��IM��F]#��#+�q�Rc��b&��uk���s`h�����5�� ��j4tuw`@�)�����h��
M���]%���i�g����,�
���E����-��@�On��GF�TU�.N���ԭw�}��Ca(�b��w������?ؿ���ӃQE��2��l�uE��Q+��W�^\\\#�d�6��9��ii|����w*ˤ�&I�s�K1�H�E�f��	��F#�@���f$��`��E^EFd���M.M!*E��i�.��:	֫0L�f�T�EB"�H�7#�4i�]#F�)K�`��B]o��i�Fjk��v������#G6]�zm``0	��cqa�z��2���Z���߿{������/f�N��>5�^8�j�:���v�p�8T�a�E��5|�������,<C��2�HO�C�]]�����Ou�P�m����I��X��'�a8�0g���v9X����c"��J��b1ϼ4 cHU�jk,��-/��^��D8�t������t(N�p0P���U����պ�J��^��i��w&��=):�!"5鏠�EU)�����*U|S�T؍�X����O\�^�.--о�n���d���FP�zY��f$�/ͤ�=^?)���빻W����	Vz9���t�f�L�Q���Y/��UjUC5��4�A�X9�H���*�s�}יI���\�eHb����!_<�E�`0IY��e���4�E^�����\���g�K��I��OI�I������2���ڪ'W(Uj�K�#���n(���fR$�k�#\jGW�LJ��L*����d�23ٜ�6HyDT�;��������,�H�i;����Rݑ���9�n4��X~8�$�B�D���p�yqw.㏷j�)�4�������������<�L$�狸bI!k��V�5cٮ\��*�.d	A@C�/~opp����J0�ݥ��s��j	��������6��C���ǹ�+�vB�п�۞���Ψ�Kk,�539���<���8����@��TQI�D������{�޹x�l6C*8�(P!觩��	?2�G�7L��^��s�u�
��V*�ff�UU�E��k�X[W{<�u��b;�l�/�u����k'�;�i�d{GK{0�ĥ7�]�s�����WQT�[�޿�?��i^J�L{o�,���+���p�n��s�&&&���̓��6��x������^g�-��G$I|��oT�׬E��w���
�1q��ߴ:-�	����67����c���nU���VT0��2ٔT#P���|�a���/��~%EV�R��ke�,�7`B��t���Aؐ!'��Ոg�<W��Mݞ�=����F���������3i`���J$���Յ�V�w���������j���-|�ih`i5�%D�����cܝx�-vr�l��H���ԯ�P,"�D��G}��,,- }&�����>�,�P-�����cǎ��x�"U��B `�m�D������P�kcG������IbD��<��~��/�|as+�q��xTj�}�`@��Ng����]^|�ٳg��wtt9~�X)�XVV�l��ҩT"��7���+��Tke��7�~�Pj�i�T�hٟ�$�J�� �T9�c�|2yW��������f��n_0���x�؉�z�!��������������#������\�c}^A�i�i%l��|C�Dk�Z�hz"������/Vk��������ew d	k�������:zzV76~�I����ٙ�^��qۍ�������n0:J%�j.���]�e�]���!��b����i���laT��,iJ	���)J������?r�ڕ�W/~0:г�:_�U[[�0��,--�v�|�氞�m`?�)׋�˛w^<9.�'��=�
n��aAWx��C��6��@:]�u�&���~���|�t8D����ߘJ��ժ0�E�XZ꼆�� 9��.�x����'�zb�V�ZiR^�������0pE�R����K�*�J[��u�dz}> �^�55}�����6 ��9��r Yp��*˒��-(ܠxz�G;�.����8�BUÕ�#�)��(4|��7����nM������o&[�@N��[H�[���q�h#>��c�&�TVdG2���(���A��7���p<!^s��;:�v��&	xf�[���ؾ��ӧO/,���0^�����o�>�KgB� �j3����ιT�^:=�]�s�++ܙ��+����fj�J�֎{{�F�l���Ս��vP���n����%�^og����O\�v9�������L��H����i��o7>��h0�@��2�9З�/��9bE���m���S�ح��Ç:t�ҥK:5*gu���+
�n����V-{��$m����mV�%�`;�Jf�a7���_WH=������t�:)b��
|�``�pJ�^�{���!+�`�/"g��]mk��ť��o\ڷo��Q� `��DWOWo_g8�y�^O 	���*�U�hb��J**$��`0�Yƕ*�b[ީ�a&b4�Ϫ��1��V,��u�j�ӳ3V�H��"A����I�Z�A_Wgۥ���?�m�J*�Սj]k����k�x�h��dy���Z��t2��˿x�����ǟd��I.I0�����ξ?1q~�^r>u�pO�kl�(B(3휩[����� ����mf�C��a������
��:��W(�<n�WQJ�J���f��˷�e{{��S��!o���	ݰ�]���ɿ��$~W�vdI�aމ�?�B���d�6��P��'�/��l�SY��u;]�kkW�\l
Ƒ������N��lIi(u��5sqy����W_-�r B����x)��$	�<��!v�m}�D�Z��B쌭�
��`� |J�3���ۡz��ݙ�m���-.gkG;m����f�ZH]�ZSݞ���-'�|�������3,��
w��$�<Y�c�N��.�aQZ����?�FY$�x���_�z��w�����>S� G����?���9�.n��r��d2߆�лX�~E�ؽ�����U��7�����}�=ۛ˳�Te�4�'|�gck��TJ�l6�فk=�DAnUeU��n�E�s�� �xF�T+����xMCP���.�������bi�U��UΖ��(�/JUJƨ���P	�kpx�������7���f�KKK�l{�1����M������"�p�^l!
��� ���QW�t���.��M��D7{��uUq"��W=n�_�JM׼>�6�Ƞ��������4|<x;o-����a&�5D0r\��b)����X�W�#�{���heG�T����ɍ���,,_��!b��G�t�z�3�kpc2_(�r�.|��/<t���Wg2���X[�c�2<{ɴ�4®��ǲH��L6�u{��~}e]��g����Uj�>�p���'�hA$�Z��
��(�
�n����W]N_0������]�ޝ�^�?����B�q�|��|�. ކY��X�n5��%�˥��	�@R,�ZQ�i���8<������8W�/��m��+F��8��4[��C�A\|�Wi��e��Sk�rU�p�5C�l�8���ҥjT+eY����|&��RO�#��'c���D	��cc�<n_�_��R�����:i���g �x�R���&�,�� �^7O@7�(~��+�]�'��F:���0w�Ƶ��u�Fd5�Jwwt>��so�>��/����?��?*r���w�옝6>2�\4��K� ��:'����h���:����9L?��L fjya�����]]]X��tW�A-\:#`�P(b3V�U��މ?��/~���Ŵm���	�X9�r�,���S�G�����A��p�"x>���c~~.��x�i���c�$ZU��eRݠ}w����ܼy��K�<�������Ǐݧ:H=� l,^�V0�X6�-F�R�q(�rz��b��̓���0�n��`�mu�ҝ.O,���f�P�'��Lٛ�=�h��+����8y�S�N�B1,���}N�/�I�Ug��DIƯ�|<^��w=;ܬi9��g����$�1%�@��J}W�u���E��Ţ"Q;`�8\��!���cm]���@Hh�m������Lʹ��:n�K�������ODyg0�qH����D�b������.��R!�7�l����fJTIT-SK&b���Fcxx8�J�}Wj��G�5�)r�O;�kmki1�������n#@<��#	WJ0qQ�S&�� 1�%Ke�~��DkBv�}�@���H4�v*�ZN2%���E��R����o��v�V@X�ok��x��z��e�b�H�X����� 	o��.��44�x�%�ڻ�I��������`Ҫ��זE��^dٍ�-LS���t�:�It�ܼ��A�4Sw9\:e���8�f �Ӿv7�E����}���d7�b����Q��\/�g?{yvv����C���S<C�G��$0\/���K� �s�� ?{�{�1��v_d�6%;����u��U�[�1�@�</�5���E�e����:X���M��&²��������������3OYԇ��[�����
| ��e���v��=G��39��f����5b4K�����-�OM&����ñ��Qd0'Y��̥���z�'?yiii��·����Y(����/O�^��W��I"�O�Og��m{�]:�@���֒l'�N��r�����̃��0l���5������)��yr}3ucjzb��v.��%�dv��u��aĉ���b:;_��7V��`��K"˰�+� ����1�l�������j�����)��Ξ>}(��ѣ<�@���ʪ�������_�}�]D^�"kpF���10)|��mb	c��y�;\�ډ�)+�7_���ɖx �ju��н��X���.���<���������q��ɱ#��� ��nݴM�	�a� � cb���59s���Kyx�Z���Kw�}�r��l��d 2&����42l�8��r���-�������mRB�3�H^Y)Z���+,�/ݞY������dC�ז�ǑJ��K��طCIĒM[D�1�:��/�k���(�j�5�ZL��MU��d�60qo��+e��\�P/����[�ϟ�7>|XT^�aT͕�M��n�����/\��s�� �xss��'p�ᢞ��%�z]c;��Օ��Ć;�N�Η���;��H.�����L����QaA����G2H��$n[(���?Ŕ���K�~�����x��*�xA���Ԣɤ���*6662M�r�ܬ�J��;�W7H�kc{mj�V{kKWG[8L���4u#�޶:��n/�� ���ws���k_{�ӧߢΕ�bZv"JU�B���}~����Z�	Q�����::����*��.��v3�w2��J�r=���--�͵�"��r��x8 6���J���
���v{[K"�ϖf�f�S�ڵ�3��~*�"̫��������A���.��n���G"���-��Z�Z��pX��OA1�G��Q�Zg'��|�������9�Z�:<bv�nM��������;y��v{����z��uY-�g+�����,�˃
�H�\ ��E�&�L)<��Z��ȯ���3���Vd��t_�,�M��Ξ���X<�3㩯�m��>�hG{���x�\�j55�z����K��E|���Z��ޒlkk��n	:B���F��uU�E K`\X+#ltadSvCeC}{z�7C��eӱx���(�<gyf�v4�Ӵ��@������W��:���wt�N�HD�ж�7}~��4����C�z���5Jh�'�<��FC�D�$� b�w��F4��Φ�'����&f[�Y�P2��H����3g�R_ϣ����~�V���6�өb[Gg���j�6���e'����vj��R��F5K��;C�
���p~QQqG� �|~���ˑ�ڮ��,�Z��1E�B������	�}'?�E�/��V��j��Pm�G�.�3��n�5��$�����9ZU��Z�e4��5uӦ�w�	g�?R�Ep15y|$5��UdJ����f7����۷o��0j�&�.T�&o�5�ǯi��nW K���t9]��\�Cb}rz�{lɠ"N�Y��X�eZ�|h��B��'=�0�R�to+�h��9����o|��/��?�s{�I�!2��i�+�b��5ʁ���8#^�)��-���}~���7u�h*�� i�R(�]2y#,*KQq�.7WÒ���|�I�E��9������J�Bk2�t�P�Y{���|����DQ��-����-���Ķ�VL\!�b��4U���Qaă:�`P�$ò�E[ƻ5�r{`���@��Iy����f*%dʥ���b_w$�,��~ȷՠ,(�5�5ݪ#	��v��PI٥�"eF`I��G�1����ZCo�&�O0�os����2�k9ť���?��?���o��3H�����,�MW{3�� �"��J\F��R��������B
)���B��n%�H	4C�cG� �����LO{o������=���9���� r���a����*�3��s�{��Qȋ��U93���X�w w��sKj�� �) U[?07�u�Ǩ�ϥ�L�,�����|�_�ªh�2���L���^�Y]�25��60�l�������o}�k_�����{�ر+�/cA�ܹsӦMء�[!� lc�7��M�����lR�8� K�^B>��Ǔ�b�d��4�im~�҅�KK�����'۵w���K0>fEqaɒ���{����_�a��u�kLM\�edgp��#�� 8h(��!�����ݍ�����X�Z�5}��\&],Wҙ�]��/��Gdٖ+�~�ue59x���r�}�ޓ�%j���Cj�n��Zķ48E�9�-�6G�1I���
P�����~��+ 
��W�^���'?�c)������^x��}��MNO�W����v᷏_��;91s��=��K$%l�pl���+"|����l4f�{�=s��dO���\�G��&�(����xP���IuK�d~�ͤK�sK��7��.뚁&�_7Q�����V&���R]��qXBC�/�<~I�X���<t!�+��р��qyົ{q%���k�^V��@�5S���\B���+U
��".��$�7�"�"��d��/[6�~뭷�8�$�i��[<���ￏ[���q,^��&įb��H����j i�E�I��l���*�b�l�^4�����-sy k����~ c 5|�č�X,655s��`2��L��ubb�j�S�6�	�
��!8LΪk!?�|�ĳ��񱐾Y�N�'X��~���]��S�(�l2	�W���8�,VV�|0teX�����G>�9f �3:%=y��%J<n�L)���Ͳ��EA��F���\�~������+�=]6����4^w�筷Z$[ow����s�=����? �2=;����X>�R!�I'eIy��{�����&��ym6�Y�B�%��d0�"T�D��˺��pBfsqq��YY�J�dr�Z��70@Z��;R����{�����Y�@�ˋ�`�ݶ3gΉ�&BҢ�3nDIE���e�Rwi�,a����b�V�J�tRF�xf�͈�m'��[�s�
�������bu����L2�����c�[�ĩ&n�����8��R)�"�)g�:�%Ň6�t5��KZT�2l��Q<SK���n� ^�kc�>�,|/Z$i�y0Q���<",!|e-�������"W��g���.��
�I�)�D5uV;"])�ikgW���h6���^�{b|����� �@��_�)��N&�q%�X�x2�F0�V��+��5:B1:5+��ᷙl�q�UQ�-��2��Z���N�ǃq�:V��p��`$���/|IUI��ܹ+��Ӊ����T��F")-*�ר᎙�B��U9f����R�%\Y.M-�M����r�T�Dѳb�D��1��j��}ێ�.a��S$�ehh3�w�^3�t�̯ba;�.�����p$(��eX�bW��j=�Ƀ���s�"u�d@����ٿ���Q�s5�Uu:�����B,�Lc���|y����(�ra�''�b�U�B���״���|~V��Ա�֔�"P�8T�Vģ��K�NTU
7W��=5f���� /E�'t�
��Е��x��=QL| �j��j����NPA���Nd��D�V�;=:�f���wPSlۊ*l f���
�r:��vt�l.�J�9APE�����%,6lD  l����b5ú�����
~J��i��S���E��&	Hڢ��^�\k�{�������Lj�������4q~^���6,�-|�LQ3��GU��>U�Y}���\�Kl���kc�P����a��������1^��9�����S�N���>���=�'B��b�c�P��w PA��is��V5:#��[��Q���<0�κ�R.O�j&��m1;fg�&��
�Զ�|x�{���.�g���Y��,�,�8p���111F5�Ա��wʥG�����؛��*>nwfc��dm��r]y��@���@F�^L-/-œ�L��P>��@����l
�[Ls�P����16��/���[�nٲ�f�B��]�K�����#��t.@1x��CI�tzmu5��3�ܶm\,L���Z}���~��������B�Yl\�S;���$�?�C-W��X6��f����!�@͔�x���'�J���9sf||~P�w`��5j�J��
%}ހ���;!*�PI�e$@����dJ�P�֦g���n8�0=��(�R���-�}�x\VR�g�gO��6t-�J���dr�Z��nX �6�۵}��=;���z��J$)ve��5!)�� �d��Z����r'�������z�s�:�X��XU�o@`K"�2x�r,��T�D"��?�����/_�8==O'��e�[<�T�"�S	��gS� |6�x�
�I1�)\��m�H�e�=�IK	z �9�ySggG��u���Y�%�4�\LX`� ��fs� t(��"��Hh��{(�4�dR�������&b��Vh���n��Ŗ�E����A4
��_]>r���m��-k��s��@�b�����!�}ǅ��A9��n`�y�c����*�R%U(�
��`���>���c�pm�J�y���\�q�������8}K��0����v���䆯���iE�,.�/���*�p����6��
T'���=����޳@k�-�!�����R���8FN�q1L�Y�,�,�\[�')�}X�G}����W�\�֪v���G���疱�9oǵ%��MO���T�}�={[����(������,����r0��;�va]�E��D]IO|׮]���z��Q�R���?VU������ˊx���)j,377���,s�+�S���]P
�(u�R�:�zG{׍7@��E#D%�Hj2�#`�a���&�s3�K����X]^�t`�����Y* #�[x�G��\�NMM��1�ĈL�`0D�;}�	����`�%	��OǪ��0+ä}]y�p1�-X�ݻ��4��ǐ�']��mm�-[6��.'�}*��u��p2���څ�Ę���-����	Dۢ,��"(�/tn&a=�VF��z'S�K��	:H����=�����>��BL�=��;93��aj��P2�z�wp�>�I�����Ç撩X��o�����hs9�X9�͈�cBq�w���+Q+�a3k��+��L;Y�0W.�~�f��*��Q�݌�2��%R��ۗ��<���̄�hii_[M��M���Up綶������]%a�,Y1�P��\�oX?J����F
_�^K������$����d,Ǉ��]���[�
)��ǧ�cx��Y^Y��lg۹sw$�s�,F,�Zf�@��FM�4�~x�Zr�z��&J},Ltaӂ�0�����p*�=��\V��"Y��qll��M�m	Pq���"�6��nu9xp�y52�n[�װ����Md+�Ba�l! �hB-qEk���gI�����2'O�ik����� ۭ�raqi;����
	��簞���������>��
x{��F�� Ł$oN���cյu�\�C�zc����и�u�F�G�Le����uCt�fF�G�h�4��Yt�v�/��/1��'B�j����s��,����1�{����G��c��P٧�!������q4T�R��%E�*�(|UMe�T��r>��.�^�zieu�f�>���l��V\�E��J���Ka/_8?��_�:x���1�k�;��8މ�xFd��7I�`41�l: ���7ԧ�4� �2L%U�lf�T�V�T�&ӽ�A�/�nk�-�b���]]-�����B���^�Wa=+�����yHUEȄcu�f@~"Q�$z]��'�D:��P
p����W/_~�7^��q�ܬ�$ˊ`���W}�0:�hk	y��@]ӳ���ķ�˚ϕ�{S�d�C7�ku���*K���c�1��l���D"�pP$�@̤EQ	���e��ՔERE 
0Ҩ�
�B*�p�Q�|
����s�B%GG՚"�X�j�n�EC������"�hf�Ak�*��#�C��-sVQ�C��f���t&%�\E�Ps���j�+�nG�r�H ��� ��"��J����5���y�	��TC�uۀ������Q�5�,SW%��vf��Vl�(���N��F�����b`�f?��On�ԛJ%{z�Xwnn	��lvv���Al x,l�H����["�e�}����g{zz0AX� 8�6�����I�&�!U�k`�E�����)��F�Y�R(�6ҹR�b���Xb�����3:v�ڵk�r|��c���x��?αjf�:����G^o)�ߐ��T��+��u����笊��M+�������/����pZ��21�M�����T��OO}�j��jy\XƸr�w�*��E���f z�09�iqƢ5+	�Ǣ�X�l'��6Jh�u``��{��E�l��t�ta�ҥ���� &���^j���U.`�´b�>���c��\Es@�miu�<��Ԝ��Z:4��dP��Ρ�+W�<��O�]���+J�6@؏}�<?Oj��P����y�TQc�����R�Q��f,<_��� �O@"�X�#�@�����'u"��2z$ �=zDC��#гS|'&&ƈ���C��rS��n�����ҡ���.ѣ��],n���!�}q��o�˒�~���-��6����pU�)!�+��L	�ĉ����"���a��lo����#��rE��0�
�\���u8L��X)Z��7ig������n����t� �Y��_x���`��6�dU�U�٤5� B ��|�3�<�,�V�V�>|mfj��{��V����X�:���m[�m��v@��%��fC������2��V�]�h� m57*��h��A�XxH�fc9�c_ð`��,�X���)�?h�,��E��G��]m�;vl�#tH��H��@��H�k���\"���犣�Gұ�_���S���4��kU��۶m��t�R�T\K�2�6	�#++K�Z�����]�h?���s�n:ˢ5�Y�(B��ɂmE����D�[RMH���$�o&�]�m���H/�,uyno���?�7t�
f��dii�C�O�:/VZ����3��;Z�zZ���io�t��T���.o�Xh� ��1MU٬[)��ё�SO�g�œ�t�Z&��G���3۷�i�2H�r@XKˋ��o?8~��݇�WcKF�,�����6��a����^S��F�����z�I�0�|6�x�8ٱ~8B-n���,H��rq9SA0�R�.�GƂn��>t"��.8��tK��_�٨A�3�a���A4,����f��G�y�f<S�/}��;q��ɓ'�ؒ�۷oЪ��  �K�;V�mC�\**�$2�7\��y�іV�F�GW���}{��}��j2˥r[�Sմ�x�����'��9}�ƍk`����~W�h�s@��mmmO>��o� ,P�&�.��xB��3�`�Q�-�"R�f������Bjeaflt�{z7mٱ}�O��|v��+����ڵc��M���`���L:Q*b�y�n��M�ӵY���k� Q��k(L�QE�����ox�W8��Q�"�)S�ި��[~��߶bdY���>K�{vmw8\R6�syo ��3?���gv,>(��M�@�V�Ch����o�cj�S��891��%!v䔬�bIM&�6R��N�Μ>{�8�7��X�Β�>7772������%k}T���^E��d�{a7��R�z(��h�F#���΢Ɲ�,�L�����8>��VW;z�g�I���U
����M��t�5�9��P�om��l�_�!%.��X�d��|��Z#�0>�%
���Y�.�h+uU�]/�,�J~��R���B��k�.xGn�q�����e�*�����lR����I+�j�d�pH�v�Zo�S��f2�N�>��r�M���l�����-[�����R��Xn�cwqE�L�S�` �a�L%�&�<}'����څK�X D%Q`�q,!�r�-�>�jx�N���V�f�SW��p�8W��P���I�(q�|��R9�4E�?��m�oˤ�@���傭�h�ȸ]��}�[�{�=��P�:��~7��U*�(���)ʽ{�~�������Ռ|D��J�e	����>;3s��qN[24���s�U�'p�����=l
�
b%	8v�޽�8/+f���B�.���@��|(�k��N`z@:\���&\	�!���1ma�����֭CCC�K�@�RYĉ��_�û���/����3���Jݺ�n�b���NNN�Q�P�Hy�'6fM�MJb0;::vlߵ}�VQ
�W wY��~q��m�Xz����<ǆE�]��!���y.A���f�z��p��S�$�J)��n+�
z�v����t�cw�!�R(y�>,,x��������s0�" �h�v�Ka��v255X�&B@���_���Sr]��.�L��yQk+ ���Ï�l@j��A�ZE�"P���-]�V�, 4�4V��KjQ)�=>��t����o�� R�bd���2!&�\��Y����-[�_�[#-��td': �,���1�(��n���������(E�mYryܲU)��C�����Y�1vPCJ����a�c�`q�����:�� �hL�8���C�S059���X,Q:b�UD͛�����->�3�@Z/�ݥ�f�0�@��EPt������(���\_Z^�G�fх��o��������������'��x�N8,�xr~%�Z6e��m�2��Ïlݼ��T,S�nߌ-�ISg!�d���)�L_�p�/~1n#�T�b��O]�Y��|��˸���uM��e�!x�î��N���i,K|��XK4�ys߶�.�d[kG��M�B��-��牟H�lh�D� _�kN�../���@��B!?���S9<GWH� �
����DE-�}s�g�]M,F"A��l�.�uz(����+Z$�"6����wt�\$��	|�k��uGj�pF�&ܷK8=g,�U��0��PU�G]�Ӛ����!��)���E�k����l$����~��/��/x�J���=^�?G"�/_^��fg�aĮ\��ySgW�?R��ʾ	Ƽ��qNdo�y!K�*�X�)QSJA=�%�X�Y��w���ؽm������:)Y79�f[�T_Z��OO9r�ؑã#�&M�,���n�+�R�n_.Ŏ��$
�g/�\��o���  5����+�B���̏�+4t?���!`���d��L|$b�N����i��wl�ݹmS4�9|�5]��m6�X�B�
�R�/Қ��k�@�Z[)MH����X��;	��Q� �)o�H��<x��7߄�JV�V��v��P��h	q��>~��j]'5[�t.�[�IS����[���?�D����b]1�nii%&����jB+؍�H�!y,���`���/�>{��T��F�چ�Ȃ��f����6��w�.-��(�����ޭVj ������z}T*+��mǿJ��\�1X�5�����r%�O���!Y�^<p��JUs9��B�ȼ�����ց#-`����@��v�®�R`R}5�=��Ո� me�0��A�p	T�Q(�n����V�T�ȯ�PC������mۊ���Ç�Vm6��g��T�
���,�}��jǏf��σ�9����y(�7S4��,�+��HQO	HW��m�����ԀX�WL5�VZ�vm����2����wʎ��{��Ww�c��̤YR�����4>��i"���=�X(��~�YP�fN	`l���z,�8����Lf>e8������\� �_��WZ�x�|��q:Z����Gvݷw�ǩ���$�����$)��1�vY��[��z���C����"˪b���L� ������	C�>�<\��p	��#9&�o��Ν������Vh�`X z�g�1_N'�V��)�'��c	iz�"�	@�-�\�w�T�{�Z�u]�ڰi��ZM��Xl���G� =�qV����.\ E�ï}��p%��-L�����qE�[x��X�v(��좲"���4��>�^.�ߴi�*a�7�|�����ƚ��/Pcŵ���gΜ���>��ёK�+�o�~?�3��Uk���� ~B<0�^���p�� [@���CjlRp!	tۨ�<�rs�C$�`��:u�)D����uww��ULֶ�[�68��m,\�O�km-��z���uut�{���痗�Z�O ,��N! I@��}��j:�H\Z�
'.�f���5�N�t��q0۾�>��V���z�3j�[*�ka�,,,,.,��dK&���,���Ձy�Do۶�	��#d,����X�x�H39��$˺*�Z-[I>�|��k#7Z�:��)L4��R�4!�*%*���펶��7'�3I!"���)���6����j�lwX�J<^��o��p�R���K�+�Kt!�F%�7�#�	��?=3.�c�n��֓(+N�.�,vJ �Xm����Ng9ѱPL��w�Px�`owok[���[�
�7(��,Uռ0���I2�jd��	FMM�=��3�pV��XW��,;΅���h4�w�0�pyy9�'t(JlD2�>������Ô��t���z�^Rl6S_����s��a��������D|��r�5S<�YXZy�b�x���.q�F�g6M�
 rۙ��d���?�`-�,-���p0ƴ���`O�=�m��9,������`ʂp�v�ƍR	Mz���4"I[�[w�Zӹ}#�Xo�1�d������(y����^�����G�P�{jǴ����A�m��yn��kRT�V8 �����w~�wz{{���_���?Ld>.4Kő3�����������j�1#��QA���%�f�m'8~J��kv�cǎ��?�P(�,�5�L[�n�[J������'Ξ={�����)_�0If�.�P��i��g{�_k|�֧����up�W�\rz@����q����@K��@�
��O�b�W���L\��ع�R�ǌEB�"#���6�[v{|fY���v��	G�[R��D2���4s�b�F�BZ� ?.��*�L����y�
��199)�ͤ3D�L�ժZ�E�������]���G6����7n]�
=S���J���߿���Y��hk�L0�F[ A0�\��a*j($��Ji=��L��j5�E����hvv�#�(��}=V���iN�H}lb�ݛ6m��H����%�V�V� H8�u,�V�4���"�]+WU�ȬὫɾU��$��t)"P1=5��/����lV�U(R�˞4��f�X����Ƨ�|����9��������y�Y@���Z��MQ�B=,�b�9t�T��UH."\�jM�%��G��T�����A�*�6lV5�>������+�}@���JY�5D"Q��TY^�J}�Ti�E�Q!��C\��'�#�)�,�>FΏ���U�,�:�;~�ƨE⤸���8q�x Uhr��No�d���5 �9���I.����<��`��%�������B]�j0�Bg�V�}Td������~��o�,ߠ'a�7��?��S����Y�ZIQ0L����-�S�̪�صW����bZlN������S3� ����PȆ�"���P8<7;���/s��g�h���m>���C��{���贀T��"�WW��K�Р���y�9�ݹ����DH�[/n����*��/ʥ|��P���"��v�Xb�T���^,� �@u#W��H`,o����>����j�B�l�UE-;�v��)��Î������ʒ���$b��>H5̩�١~���x����ȵ_x�Yx'X��.��X0b���=����[���mإ��F�tS���0��������XKW�t��p���/eS�	UcLjUʫ�rD].��o��6K1Uf����F���{ ]Tp�����������s�`#���t�r�L2G\pz����y�9���z��XL��(V�Bᤊ�K��<>ܛ� F���$"�6N��{�}���8C��$�uQv��q��q�J�D�۰��l��5 ����b�����a�r�-�ɚ�׭�^]�t;��&��*@�<���019�ʫ��ܵ�̫5Z�Z�Blu����9������w�	�I�0�X�&��2I�Ø���r�]�*e�T��,�S������Ϯ���GQ�mY����V�Kf��������>�eCA�Jȴ(�{�ĽP���$d{�����x<�K�.�˒�	�g���=ݽn����Nn1cًn�$^:;����eX?*͉�5�`8������;�y���/���_/c�GU�<n7��"1��\!lcM��zz�&�?�	���)�$�]>,��Ņ��W�psT6)d-D�Z��aI8�J	���;w��C{lP-�^�P�T���hA�l~�7��I����3RVk�`0v\�><55��)�.mm��c��~/X_�X�;����f�1^Y^[Z\M�s���h�Tg�C-VE:����]$�wEN��!���H�(�DIܮgCq�Gƅ��Pď���?�|��%oa^��/[{�#�Ν��|��W��{��G�W�M�"�5�♙�%�ࡖ�3�Ss�36'�IsJ9w�ơX'�����D��P���.�Y�S^'��J����S�����9~�"}���=�0�Z��:����Q��a�|��O~�a"�eB�z#(>�nRCטc��AP�)[��2p��V�A��RΕK���bbuff�zWWOgGowwOwW/<�������|��^I�:\B�O��#>��tz�^�[��b�Fp.6!ss�ϟ���Cׯ_�����?�� �Q,f�����-��}E~����D�Tf�����T&j�E�-�.U��	��U�M\�)���4:D��}"�Lq=�!P#�U�uU�8ܮ�f��&���_�����i"����NV7A-��&��Xrm5c��&�N�t�&+@#�X`@l�H ��Juv��"!uq,i/�牳v��Uq��`8T(m���>78x����f�٭�\��L�6Q瓩��:-���Z�����?��hO[%J��hii)�T�b,�T2M-���F�hD؀FTw�c��E�GQ�Dzn�1�l��߆����g�GcC�-aٴd*y�ر���O}��ء�t�˟�Ӛ�W|>ﺆ���i����*@���.x�>�E"���ӷ���H-4�֨O���7^}���X��r��e�Ԥ��`[(�pꩧ�̑N�@���6�NO�Jq�0�N�x%uY�P���JV��̓��tN�V+k��T:�K�+���j߾}##�vqR��ڠ�F�<�9�1��Ν;w��� �.V�ݩ���A#��;�n����^�~S��Y��;r��k�򅼪bP�	Pf������HB+U��g&3 ��'�>�.��׾��n۶-_���|�Kq���\N�C�>�J鈀L������xd�а��X�vKk�R�\[6{�v����Ea����3i�ℴ�&���O����n�d_:���������kR�I@�0�33s�JV���w4??�iQdҍ���B0p.�<|���N����ь�!\�59r�̹��L�A�e��H�s�<j���p� �|"��9<.�@t���3�;�z�B��lrU�b��qo��{s%�F"g�NL�`N�K�3�'ӛ�W�$`]a��}�vG&�&�k� j��ͮ��2��o��H�ht��JɕJf.\��~�	]68�Y	�W9{���c==}���QP�Ӏ�$�]NgM�z~�(��m�Z*c���H9]h	ұ9I}�A�ay,>+w�H�ʺ�`��O���"�)DS	&ϊl�'u�j����O>��/��x%x]�R/�s@��f��N�Ϥ�~�ar(��C�!=�� 6H�شOkz8�j%�E�:S�V�\��aZ����2�a"a �(�������k�]]e��Y7�$�lhxus�Z�
���������{\*�����Q��GHVY�`Q�S����.��P�;eM�P�	��ġC���{�}�����+��Qs�O�*1X$��Ѯ.J�����9�%�C�
��Sc찐�Z�@I6��PWVW��(��F�!!1>:��l�z=�L&u���O��>_���*+Q���J�bU�*�C�&��,/S/l7uͲ �z<��=���i��Xf��IA��M$c����jf���x�Z3�O�\�z��EٕnT�Pڨ�'�BI�j��x���X-�x`��ք����梾��5�ϰv���T��,٬� �!uC�?�\���e8; �������W���iaUXTy���t�V9ύ2���R��X����G���C�+n�ɺ��Fpl+h����-
���"�b��.�����.]�7qm�: O�T�H$0^.kB�F$�T�;Wn��$��cm��a*���/<��C�VT�����>�����~\�8^ׄ�К<��.}�o8�c��������^�Jē�3S3�s�Ks3��t*�������NeH�\&�T)W���W ��ѶP�Et����/���^�>r���W^y��g�}��zwjj�\�4����22i�2���C����>!��`��3]Eh�jZ��_-&x��p�������
�1���ry���H����X�]!i/��a�bw�UR�����n����K6'��b3�u������ѱQn��9�,�H��OnL�eZ���p$�?��%�Z.��J�J��j��`Y(=�
��U*��.��
 _��n�ՀM���?$�KUz��@����o�:uF $ֵ��(I6��
�].1D�?�QY�$��Ñ��˲X���9�` �!�B���M߆��O`/�LF�$d+����fr--�@0��k���g�s�� �]�=���"=p�.�[�^���{q�IN��bxDɍ
F��@��]�HX�c�m-�������X&���]��R�K�F�������x�ĝ�����a�!��1V�8�Ewtvl��k.��L>�IP����'_���>������4LJ$����..,./-��b�*KrgG��fw�h:\���?���Kq�`$5_so�:�z���������0w{����� W,W�&V����R�n�n�O��t��U5����݋� �Ϥ�϶��������?g��.���n8dXo�h��h�F}�1��J��ej�,.��j�]VTWg�V��2���*��6[8�D�a�E�a�h�*�*�`0�k�D���W^�ɾ��������w�Y����F�Ȓ/��{7mڼe��"�RPȦ�t��_B�_�T�w��a��5���hk�P\Z\�7��@wG.,f��r�C�/�㷿=r}d=�Jl6 
���G8�����x"	��ȉ�r�X2Uq�,|"�������AoPQ�>���r[6P��V7+�j����C�c@��Z�������?6��>fd���ը1}�d@����
u��
|V.U�II�'�
҅qƏ�p��)����hd��e��[4�דΤ�Tf�[����~��cǎqx�(�]_Ϻ��K�e1Űj��O|�05,l�U|LWDKSI�i�Ev:��%�7�tN���r<nl,�,)N���`hV;L�]h�?~�����-/-�w7o%*Ϩk�l��Ɍp�*wx�'�a��X.�*f��p(�. ���Bju��Y�
#�P>��m ����!�X�R�t(�w��2L�+W.����w�~��3���s�R sdK$��|ᓟ�����U�"��5�����$��\6e�xtM�*��U������Vc�B��uiz�h������P���������WNR���Z�|C#�D�3Ҭ�)`ѪZ��g>)�&�;��6j�d�a�Yt�20�(f�8WG��8�n�`�I �
G0A�E�(���Ǐ��ry(�X�zSژސ;�I+k�
�y�`(R�$Y4U#f+Sx���e�j�ͭV:|�g�q�"� �9�ʀ�G��`��J�d1
�t:����!�o�c�O��ĕ��VMM�Z�j}�ݳs75gq�����ɽ^8S7LL����=�Ӫf����i��S��Yn��7�_�/��{:��!+��1T82e�
�o���z	����3CCW1��/�� �2�%�lr��{݁p����������Z�ۣmm�h4�"���ͽ}��m�����.����I�bsj:�<�4ɠ�/-/�,�^�|�ҩ�'�;v�����%�9��Z�$�z��1�k�)C��+�J֋^[[���?�sVj�!��������p8̹ݜ'j��߶,�֩m.W�e�6�l�J6�[YY]XX�������~�ڵk�###333�K�������S㰞���'�;��o������k�8p Nbbb6���
~Kb�]���B��Ù�HD;�1M�isQN�p���Iňڟ�ס3��B�!��%�'w�?Įk0KTv��E��ӧOs��KnA���5���'*$�)����VJ�bJe(�"�@{��n,��b�����ଆ��������3�<æ�.�& ��To����T�NB4��͢��R��L����x�xp��0�5������� o�ڌ9r����>'���ܺ��݃ƽ>@��0`��z%
��)���NԴ�5Z.�$*�0��T���&s����Z�mۺ���{/�olkm��w��o�>�{a�	���}q�0#"r��۬���>�gna>�'ڀ�����n��E�,�+=�Q���W�\Y^^��!>�
��}?{v���sss\��I䑿�]�CK�-��a�m۶�K"M)`k��3�Ɓ껂A��#�.H]�Tt�I��U&(�Ҵz{/\���o|����|���wi�rx�����Z�5�m�V�̵�U:U�\����Q!��z��n��V�:�rR:�"�q/6����@�|>�ŋ�����kpp�$ �%gjw��@��t�S_ow���b�\nok�\�j�����|������Υ8,*������v��|>�H�H���}fv�?�с�Tg���ހ!��<���{"�:�f�ݝ��X� lO��0XB�H.u��ħ�\9��s8k*p[ޝzE[jU��W_�����$�$å��u�?����ڵ�٘Y�-��R!VBM�"����B��x�8�F@k��b�
��jmm��y����.�-�wf��qwx�O�1W�q�����vF!���cĚ0�x�4+�R�Ӊ��y=�RW�����/���{������dW�~^4(}��;�U�ج���O.W�k�f�mH��޳6R]�Rg0僀~�G�h��m!�������D��=R4,9��L�Y"yhMh����V�u��T҆uQ�/U�5 �T&������.'l<�?��P��n��[�������z�y�6�m����d�J�G��G~TP0�क़&����/q�n ���"�=XL!%鐨*�D����Z�i�,ˋ[���?{��'���Vk�ێ�!%�F�`o����\�<i�h���0�t�_�HB���)�.�8#\<���7Zh�hp-0��_��S��׮\�K+�������jݨ�3�%�v!	�沋;2$�-dԛ��wF}u����KN�/����m�H͙�L~jd��7w֌�ƣ�K��СC�N�A�-۩�����h��N��Sj�ۣ��� ^�h$����Wn��'~k�Ob��L6711y��ٓ�O�<�v�̙�33��r�D�&��b�,����؏\,�n���S(l ^��������yN�%B�m�2�(+�`��;a�D��>>4��can�՜���9%�w��	����/��9�>F���CCWΝ;����|�������@9B��̞�����ZX� B���%���4�z��vP{GJ�6����jUTIB���n��������j���a1[�;'''���s�4N�3�0s��� ��$��p�VE�^*��T�\����c�&&Dx���ZUx�$d �oD�ώ��v �����e!)#�q{���x�������xVK4'!��L2���M׎5KGH�I`�0��U��u+@������b$1�N2_N�݁]��s��0�傊flmЦ�IGIk�|�i(p{�t�<��Re?�p�4��Quxݺ��!^^ZNg�===�$�i�gjo� 3 |�������U<CrҲ|w��d�<35�J%�.\�B��,���K2QN`��J�].��,��,,,Ҙh:\�����F���[V����߂'I�|Th2���]2���i����~)uU���Ӛ�鴔�|w �5Ғ.HB�������"
��DGG�������^�%WQ߅��,a#,-/�~D[[�Y ��gt�/�v��i�MT���%��a 4G�1Px�P���b����a;\�:�_��>q�$���lVέ��LMM�P�D[[[Z<7�<���^�� i.��J�A�R��7������#�(��_0��ѵ����˿�e����.8��`*����XE�޻�@7�`�Hu�d'AuQ}�����[[XZ�U)�@����p�%�
�/����������tl�t=�U=^Kq!҉V+�?�8M�$��`	qSZQ8T��̸�u����snj�Hѭ�JBI�����Dkr7����=���/��������%|�Oڲe+x&�c�5����P.�]�Ĺ����Q�#d^�f�+�{����lJt�W���c?�я�y�L&�뷉~@�Ǉ�	�<�'��� �`,^�S�&�뺩"X5
Q&�*���P�Ę���6'#UK�r�r�������Ξ���+�1fD0� ������[wn�4!�M�q|e&۬����-!������z��b�J��R�.��'fL����[�60�d*p���N͌9�v#��0�b�׹��C3++���;v��oV�5�j��uA����ƍ!Lf�lS�tM`D���?�4[dr
TM���|��A��<x��D2�ue�>����m�b���n�=��ޠ���Ȥ�R�d��\���K�?�a*��f��P�������&�iY�y}
yR,x���꙳�pa B�L�f#Ln27�t"L*3�a`DyySJs!l/�+�24�����F�7Џ�o��lx��q۳�W�����s��s� ,*`pE�Ul
x�0,��h��K�.	U��ɳ��N.���?űI�֕��t,-����_:W��������������9q��{'���~mhjj�T�)�Cd��{MSô�kYY���r9 f���p�������������q"�pXKKlP)vGy�����̋��1�XD�)j.���`j;TJc� ���,u���*�lfee5�STI8�z�)�� ��?�n���_f�H"uU�<��������v��&�S&�	���U�xl�N0�uq�c�t9'�{#%�3W(>���`A���7�H�,��X�9�	SK��~V`6  c<�(��"LZ�z-'��B�:�`������6mz�W���ob�r��C�w9�VdUWH5����	~4��98:���:� n��< �qO������D��j��^Q�<��~����a�����Fo0�M�����7����۩x�B�>p&�Y��f9�w���f7%�C��k��u��
�f��遅=t�X�2K>���+�y�P�@/^YY��.iok�9�qN�@I]�|��gU��C0�����pwuuG"`a��;��M��˗�uE)��wr<շ�y��4����OIY�~p0��!��g��j4-��V�o�#,��EM�:44�o|c���� �����]��6v��������z���F)"�(n�X�	W�b�8:p�d|�� ad��O��}>���� �_{�u�*�D:�i�u�z�<>L#��FWVV�zz6Kt�6k�����\���` �0�p�s�ŉ�]��`^(H9�
��oO�۷/�LQ�Y��-��1Ȇ��~�a�Ν���Y�T��ǘ�b��u��a�oP��,Z���F(�!��^E��A�����;�����A��V�5��jG�|҂�����1ٻwo  ��j�9V�b� ��
j�=�����P@Yj�I��` h���*��;����ҥ˜�v�J.��� ˅_�x���##dW��^�	���h�J�S�$�38�ѵ��,�y��_�Ű�����]N����J#H�E;����͛7o�ԇ�TR�Uʮr�Hj��g��玴B�R�+xc,H`�"Ӡ9]�T,�g����n�U`s��
�����恎�N,�2�u�����]�(IZә�P-�ق� /�'�<�����"���tY��S����g�������>?q 6��^�bX�hE X������;��6b�4r�i��
,�Vl�ZA��sn���SҘ$;�\��^��݆���,����ٹY*�6��X�>�fV��=>�������+`YF���R����;��p�Xaf���4]t��*���d2}mx����X��D���%�tQ2<�g;0PV��e�ce�a�񡗝Oԫb#��n�7���2cn=`�˙ϭ��[_�����֡��F-�$�s����7.7=��.,��,��	\}*�0uN���:?x�~e��ȍ���L6��2�pV�H� �
���%�p�v-�+�V�_��|i����9t�ĉ�/^�H��e��L�/��B�L� �-r)]L~�Α3_����YV�������}���@����{���5��cX9��L�~y.d�PC�#O.��ڻ��$����{��)[���\���h
�֟ߖO�o-���ߥl����Ie�9�-��I��֩Z�a'����"�.H]�n����V$_�����'a�A�^O"�|�����@NFp�K��YAN)�X��L"Og��-����C��Q�Þ+�����x�$�K)"5涧�W�d�0����_<�̳ ��������]�V7���)\Mh�
[�U��}�8��Q=X!�Î-��B����jԝJ�!��twwwvv�M�>�ֿ=�C�+"���J��CCxWZb�5p!x�p8���y`����b3��ĕ�3�JUu����'ؙ�{'�u4��^&#p��[��ַ'&&X���A�����j�a��Rq/�DF<
6����{�X��ZI��!bW�GL(�I{GgWwO0^\Z~���?�ɾs���F]#A��V��.��UR�2F����n���+ ��l&����E��7�m8����X-��-��]{��c1#ֿ8��Ϝ9�7�7��;�"5��53�[�V��JWggg���2�����|tH�1t� ����e���i����j ��
�:w�,��[o��jFU1���Z�f�m!i�������l�%�e` �L��V�h9�w��^M���
~7'�#�\�`�� .��塧����=�r����.P���q�Jra�ɀ��x��h�4�݆��s�I���LX��3����t7�~)6��ӑL%���;߾v���Ȣ��v �����rՑ� �;w��� �%�&^cIn�W*��fs�K���nU��Y�#�~��>w�ܿ��=z�[H}8qQ�@��qT���aKb�ڵ���F��	>���|*�,�E���6�j:�X���D(Q�N�B�67���sσ����=Uk�f,hpi#�������۶m=�g���t� ���a��Y)�*����I0�Z�)�˛�:�ٳg��'��dAa�v�&���X�����Ľ����ށ�����*���sM���kEh��d��ul@� �Q�r���9�k���N>��G��G����&B��H.����9���ji1��֭���`�~�c1+�p�������	���
)I��D"u�¥7�<p��{�;N���ǤX
�s�88��������M}vl�n|���h�fa���h���6S���$���
󸰼�K�E��Օص��W�\n�$�w�)/Jv��C�
�&N�8g\'�NQk?U���$:���a�r�6m��φ�������Z�Ӝ��y���9�LoX3�`����p�[��`���
����g�S�����������W��:}��;t��ो�`<�g�����(�gl���Еk�W/�?q�8\ƩS'��ޑ��J^ğ`�r�,�;�_]�
�@���[�~T����7Nkd
Ŀ������_��_��_�F`�݈��=�䓻w��L��E&�&Gb~�CV����?��m+�NrB�hdE�ֆ�(���0:����+|�f���R�__f��r�X]D�)`/Z.�u���N2qN�+UU
=Y���!�-����*�XD��/���/���K/�����_&m�aAYX�*�[%
t���ut J����/�����=�ΎhKǢ6o�N5���>�췾�-�y>�K��]��fʺ�H���Ak��
�b&��O�z��ܠ�fxz�1��8R�\�jw:�>?@@0 ���瞽===7n�x���^y���x�c��٬�ܵ�F7�4����M�%��I�S�T\�m$��.V�
%{8`���|���M];��9������$izz��W^y��^6U��tYz���%��7��Z�ff��c �D�,#��UqP�%'�y��ήΖh[K4�����ա���������(L-;��\&�Xw$�����2C�u@�r��E�Vs�P��')w+ դ5'�k��-�!�B���W~$o��6�'�����p\Ɋ&��Ņb���p�A6�"E�T*�RѝąUX<�@�MGyN�X,2`}��q*@r�C ���n������������,V���	vi|�Z�1�:�[�:�z�4X�P(��������~��9z��zǆ�5�f�	�b�@���ٹ\6p��ڎ��GY:�s�2��X<K�C�-�*�:��._��o��0S���� L���w<�4�ߙi3ނ���`��������X,��[�Tu���d����$a
6O2q��8�}�p¢�~b��y�'N���-~�C5BM�+n>	��#�s�N.�=�%q�/��pĒH�1�`��G2�����9؜����3�=w���z��n�]�&BF_�	��hg2�K�����'ħ3�b�\�T0܄� �)�M�	IRE�F�`���`2QOLN?q��^|睷9�Y�B�>�Q���B<�=7u��/�� qmG�Bc���(WE��t�Hb��a9�ӱ��-_|��=X��|>g��U�7�r3�6����6V����X��O�3~���o���w
J .cK�G�a>�����f[�.���P(d'&��=z��[7Fo4�rk�;!6��������nXtn&S�
�����a��tjz�»/,-��x�VCa<S(���� �O�:344����59>>��Y�0��F�1�'kuss^��8I���)���ƨ2�0�3���߇_�|��Y.�0^l_X��<c�Po��J���x�H	k�
c@Q�ud��4�)����7����a�·�r�B���P� RA:�Z�_�~���k�.]���̙ӧN�:q��9|s���3������^�|��Е�Cs󳢷g�
��5z(	�ibe�`�A��TI�"�'Ycȷ�Am�J���~x[��O<����:�$B��}������s.���.d^��7׮��4pcJ҉���d��:�uŌFc���S�W�S@񷏏�Yx-k�$��$�qg2��
y�T2�H$�V��T���IQ8_(��d27 ���-�VW�Ξ=���_��x1�9͉wGKL�(i]�粹t&].��,�22@L��&�K,j�I��p��T)Op:��������^{���8�G]�E�݉�b�#KC}^3������qܯZU��r��/�J�d�b�������*�E5��t
Q�F�����cǎ=���Ǐ����hC���V7s��ܖ�$��eq@9x�+k@��4�RŐ�\�k|�)w�յ�fP�*�*�����/�D�unnv�5�1#�yG�H@��Y	f�8�ύ���_&��k*_,b�s�+�[j�O/��l6���� s~��wT3M��Fi����^��E��ع������UQ��j�.�����CA�5 �_&P^ħЌ�O��'�����"��C�V5�_F���mG���D��aǭcy,-/��UHj�G�Jc���R{(_HS��,��C�.�������y�����:x
M>E4굚��d�a������SS����VV�x��qe9��VH�;bs��M0�װ���@�H_4��%O�o"lqM��8̅���dR��J`}�,�qy`� �?�� �����A��9���|~iii�����Q�ߛ��Y��<>>���4�qYb��9|^�N�0��Ry]��`u�RZ(C�rcd����ǎ��
�b�em�2�AH ����/\����8`��	l���
�1�#}�ӥ`Ə?������7''�8�[���r�f��/R�}ff���--�`�"d�1�&�8�zt\f�E��* 2	+c4�����7�<�����1����p+k���0���$��"lkk۱c8��a������D�Y$�Q*%��E[�#v平� �:�?�Hĝ.�+e����i��< �dAQ�X(sx�*1g����vae�S���!
��_U��bj5'B�����ӧϜ:y&�V�	Hm�8�.5T�Щn�eh�tL�V��]˓U�ϛ�֭U�@�‶<���P	7��`��Ј�f�b�C,ĕ{�j��:-mk��:��lP
y������#�;�����s2�V52����7��9������}F����u��ۭ�	�&�/��:sdfZ��p@~h�/_������֭���?yB�����#�����ыW�^v��k.��5Ew�5q-[�<\������&���l(f�=��ܴ�iH�{�H~;D�=00�u1\�K�^_���ݭ����:z�Zw�9��B:����0��y ��9�d�W��ʟ�{�d��Dt���1�cׯ]1x�_�p"3�n��fn`J��{��"��6m٦~o!�_1��|m��Q�j}y*kaс�W�ąv@{r�"9�l���o���[�?���k�N�������{����[D	u(���Z5�W	?��L�%��93�Ep��gqX$8,�5�tݵ�DP`����FF�ݏ���\>�}�\�k߷Mt�d7�Ƀ��~��~��2@gtE�BL�X<bȎ
`�7���� �ΊN��e���;Y���/k֬i��i�n4�$c�˭5�t���ԩS���AxX�d���lw�"1DܺHK���އ��~N��Z�V�����D@�#E�[���/k�֭[����8q���͗�LM�2���a�6.�ԒF��	���ٯ.���-�r]|�����A�$�ʉ��׸ڪe+�[�N���#G.\� ?�O�k���u�\aNT8 ��io�����u��]WB=���.�"EQ�W�|�ȩ��_�t�;�z���zk@��1����LDTx#y�l�t˹�6���;�|jӦM�V�i����l����u#t.��Swܔ�[�}��P2Q��"W���⬞3(-�\ꋺ�v��Ȭ��Gy��'~���b���4���K0��`���̩������3x/��̜����0�)��A�m۶�ڵ��GE^�=<$�x�70D��?�̙3g��0�zy7���=�°�ʟf����"��1�K|J���o_z����=��CH�z�|���˺���&ܾ=!�y��B9�>��O?1v!��V�0A������?���ݻw?��s�>�첑aag1������[�Jd��/@��/���s���������O�>����&���%,X��3��d3?�_����/��QV��¦[�L��:d��@~������񋯿�ZpQ�w�vr����;��A� r=t�98oܸ�����x����T{�>�A�c�{��u���:���?����S�n�������*[�o������o۷oA����j!�p��P�%�s�ĉ3��8��7�.\�bD�sr��0l6�Da.^=��\��)Myn��|�ˆEC��⋯��ʃ>�jժ�(.ٻu��d��3�j���uz�qS8],p9��'�G��ؘ��#/�P��8H��L�!�9T $d�Q��o��v����3ψؑ�z�
#l��r���S�Zg!{�����w��=&�5�U���\n��F_m�u���R���}0��b�e��&���./(�!��G��2�߇`�&.^g+d"�(����kG?��M�C���h��[;��Y���SnKRt`C��h ]��7�] ��u}C����G��&@����Ky���(�J=�P�<MW�_)�u�T�M|���X�bDV�؎K���:�s���8�޸&�7o��������+��j'�!���og@��vu�%��0��Z��$�
�N�9��i�/X��,�5+r{����O31Ŭ3|_]�l�7�j��������4`
�ї�Y�y���GäI���^V�7'Q]��h���`6�E�l���l�)fUc����A�sSG�\�,qeo��W�k�*�Ŏ���%�n;�����
���)�f�h��Mg�
ߠvD�r�՚.#D�9|�3@�·됞���x�tfV��'\���MEGJUvu���ߎ����򈊖��Lc���ؙ݊oq���)�����k{b�Z=1u�^�e[�$B���$W�\(�����J�,�(*�L�UKT�����ש�A$pL��À�P��g׋�4��=�\�rݺubE�8�&��S/[��ܹq�X��?�;w��� �L/�`�ov+"?�ܾ}��Ϳ)�}$<�C��쏘L���h�������Ղڋ�~�F���?,��Ν;�lH��hg�弎;&��`Y�6ͪ�WCnBu(̏�7V޴i���?/�"��B�B�ρ<Q��ɓ'ϝ;w��w��C=�R���,o't��O�ٳG�,�R�ͻT�eK��C�n���Ϸ�����v�n׷�I�z�/�ۚ���8P�r�:x���7o��ٵkװ�a��%�ٸNV�R���/���������#��Y�Ǎ���(��]�A�x���]
���"��弄x�6s��R�;�7A��NT���h��������,���` �ȓ�u�i�͢����V��<>��AW+���T��3��b��1����� ����4��t�w� ���x(Q�Z��\	a�K����s�M�Z���Vg�v��B^"bGhf����1_xᅏ>��HtZ(�x�����н��r�0��r1�S�-����8�	�G��3F����y���MB�n�Be����c��"�f��{U�-_L�b~��ա�0��w=��h:�G�����J����v�4ej�Z�Y��5�}� �pm_�&���ҔO�^y�;oUj�6���J����@�B��A�j�=�^�n3�h�^�u�t^��%@�(�X%Q0]dCR/#�����
O�3����~j5 k����aE�^4r�����7�_x|����!CB����S �&%��dQۜz�r� /5Z�0�~`���Z�`���������������~�Ș�I,S*>9­+W.����5%�,]���������o`��8w�����%ws��G��� >���$�[�� I~#����鐩����}����d�J����B^��KhM��N6G� l�F��!T`�n�'X�ŋy�ȉ�����߲e,�!����B�e�����]�r�ʝ��+�M�Y��̬[����2W��/�M��9�y���ڵk���QR�N�S~ܐ,l���{��Z9��G��Y�O��]�<;��wB~L�z٢�72�K��iQ###X����|���k�I?�I�����lW��5�i rA34���¼2#��jZ�kA�vg�!��� =�Ƈ�ݥ�o�g��ߤ�q�y�4�tL�g�љ5�\�Z����9��f����Zu� M��z��Us���LR4���z�#�'�:��X�����O?����Kl������'BӐ��	�Ć�d�G6��?�{AK�<��g�`��1aĦ4���mb�!���1�*̏jO|x��� ����Z(��̯p��רu�1Tz$��nST�Ŕ����FaEr�U�<�r�� X��+�QY�5)�"t���ι_t�34��u�q�l`U=��W��K�ѭ3#B��R�����n֊��N��7����p��$c��0�Gg;��k�ȼ|��y�ݠn#��͒Nt�Y�:	#ϡt�h�N7q2�i���~�H����ف�~1	rQ�Nw��Q�b�
�5�)?�����g�~�V�e���qr�9�O�zm``OT�9kb!0�t/X&�ئ��E�X�����g�0 ��L��2�1�!DPA���jF�,�ȱ�4R��y��hg��R�d3 ����]�T-����@:%Y�ǝ)g){��*����ҡ�`Gρ�_>��B��,X>y���Ɏ���1Ҩ}���;~�ΐ2�1�%L� ��%�@ �l������rH���?�+:��-�$V+a$viB�]-��G����M�;��j��0Z����D�Ү�_V�"2��pY�}�J������A�y��v�E�J�E������o߾-�<��;��ݻ7�7�E>��o��`�5�4�#BF�{�n��P4�)���-LؠA_v�z�Q���f�3j�W����AUF���h�/A��1�hx�"�ӣ8(�їi�7���"f��q�j�]�ځ�(E7�4:ˈ�}�.�Վ��t}�a���31c�Nz���85�)e|�q;W��J��	��(D�6͆z3�	�0������#y���ÈV�v��ؗ��$�8/Σ�XMǎ����cQ�p�ҨG���da�#=|Ʃ���!_�uZ��I�0��-�b^Mj���wR���:�x�0қI&Q��*R����BQM�h��0*P��x����7�?E6l� :��Q��as�0Ð��Q��9ʊn�tل���D�p[D9��83��xͧk�����}��Hb�i}1Ȁ �P��|���{}�E6|�or�w�J�20j���a���:C���J�ח�O��4J)^��=�Q�$ ,����zcL+�-Dغ_6!ӅٛQ�&V��Uw�"S�]�uюN-3�S�4K?T���~�fNQ4"m2�{L/
�K;��PXTZRc��I��hMF�5�BnD�r�#��cm��WD�* ���4~�q@S�5kָ?��/_���߿߾}�=s->�jll�/����O:4::�}_�z�|���^yŊi��_�Mm��ƀ��6T��G��!�3�\G��I��n3O%�+J)AʔPH�f��Ї =�l���h'f�A2�L��^�S�{�z-�1c�V��+s�S�^�l�}8�&��I��jk��N��R&��**���픨����S��V(���9�`+L Q?E�zSs�k�L��$Uj�*����Q�q|�9rQ�{�����~PN�TP�^ሹ[�@�J�Q��������e�@Y�:�g��u��(����� e���F@��
+J �A2�@���Gaf��Ui�7/Y������7�"cB{*RנU�(q�y�պ�����IXtIe-L��MM����i�gzIHa�^����T��kM]䗨o+�9s㴖NB�Mu��|*����oB���gd!�3P������������5e �oQ�����+��ƍrj[�n}��^���^����9�����.�O�5���%���H,�=j&���>Q��3�¨�x�nYF��N�4�Ja19���$)m��:7"ш�j����'��5K�vA)�iծ�ݠ��ƌNu z0��"��Q#Rv�e�ӨP��GN�%�LZ^� N�fƐ�vV��^{Ԍ��t�۹��p&i�䇄5�3���T����J����L�!s��I�*T8�-.����cc�b�*v�1�b�>��|ts�zX\�v xf��]�kz�B2����:�H/�,SȈJ�|��L׆n�%�TG�T;���w�
y�$B��L����@�0��7Mo��m�v���Xkn�](b�|DTJ���hϰmz^t�v)�?��N��EQ�N�3���H��2�[�7J�IиSǎ���2l�-�u�V�x)��3�Kk
6�0�<)
�X[z�Mce�G{ZUñ�N@U���ũB��$�v���5捩cIϦ,8�k�.k4�)´Hu���	j���H�^�E�c��LD��B�3Q՛ZbG�%As�Nߋ�KM�h�OgW:����0s�x�~E��^'���N;��m�kZ�3޽{�޽{��ٓ�c�]3�>|�ر���K�.�h���l0������)���1`�g��&8劕��I~E^x[���cH�ϣ������Q����Qi��`��`$�y$X�{��Y+���vcҟ�@6��1�AGQqdeݥ0�-��L.�I��5�K�2ث2,Xe�@�Jh��u*Q2�@+:ׅ�F��6�ʐ��Fl�M����-��>�Ϙ���Q���!��`ZS�0�A?˸MB���.���#�[��;���������Z�`�3���\���S e_�>#����)E�Lė�:��0E��L3 �R��7�9�!�g��V� ��L�Ma@65�1��~#c�iD:�®G|�!�!&0%�Nh:�`�� ��"�fZj�I9�SL)[4#T$D=���v�o^�P�,K_���+�1�3Y)���aA�!�n��T�v�d[d�S������~=O���s�
�C&�C��no�0�Ͱlav���uAW��8򬬝�+f�򧑔�G!�_���&1����S�yMSګ��B�Rܑ>u�V^,��R��5�4
�Q�D�#���a�|����lK�c��LP�0)О�(_�����������]�M0�ei�U�}M��t�1�LK���sϗ/_n�D���uB��_�tB�fpHZG��MD/k�7	G�f��Ka| �C}�<�8G��O#��t�SӳN�p������L֨>�B��h�A�zx�ME߱cǯ�)���
�֮]��t-]K�ҵt-]K�ҵt-]K����_8;�y�ѱ    IEND�B`�PK   �[^W�/��  �     jsons/user_defined.json��Mo�0@�J�sl��G�܆ez�P��iב;��I�� ��4́>x}1,���IG1#6b
��؛�:�+���`{��,�R��0=�� 6ߏ����S��p�dU݀L>bfS�����{�}��V��1_�R7�N�¨���N�Ґ@Y㫭s��Ė.���O歉�	���x���ܝm���=b�`ݭk{�9
7=mm����p�B�i��i�ؗ�9�@��k�5���5a�v?z�|\���;�d;)
Hu�s�(�R@�lx皟����\����
qZ�Á������$􊑞���^�b������Cƈ_S<0��KF�����WX"�b>U8�*-pZT[�����i.Pu������ܒN������5�:����
���3�f|�W��>c���x��ѩ������`�<�3�+��rf{�3U�������L��|�x�O�'��`�h_.�"���/����PK   �[^Wu����  ��             ��    cirkitFile.jsonPK   �[^W���[�� f� /           ��  images/8959c7fa-44e8-4699-8891-15a891fa383e.pngPK   �[^W�/��  �             ��� jsons/user_defined.jsonPK      �   �   